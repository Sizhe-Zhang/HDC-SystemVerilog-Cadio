module hamming_distance_block(
	textVector,
	computeAngle,
    index, distance, bestMatchID, argmax, done,
	clk, rst
);
parameter N = 10000;
parameter PRECISION = $clog2 (N);
parameter NUMLANG = 10;
parameter LOG_NUMLANG = $clog2 (NUMLANG);
parameter INIT_ST = 0, CNT_ST = 1, DON_ST = 2;
parameter NUMLANG_MINES_1 = NUMLANG - 1;

input [N-1 : 0] textVector;
input computeAngle;
input [PRECISION-1 : 0] index;
input argmax;
output reg [PRECISION-1 : 0] distance;
output reg [LOG_NUMLANG-1 : 0] bestMatchID;
output reg done;
input clk;
input rst;

wire [PRECISION-1 : 0] distances [NUMLANG-1 : 0];
genvar i;

reg [LOG_NUMLANG-1 : 0] j;
reg [N-1 : 0] langVectorsMem [NUMLANG-1 : 0];

wire rstCosElement = ~computeAngle & rst;
generate
	for (i = 0; i < NUMLANG; i = i + 1) begin: GEN
		hamming_distance_element #(N, PRECISION) HD_element_i(
		.langVector (langVectorsMem[i]),
		.textVector (textVector),
		.distance (distances[i]),
		.index (index),
		.enable(~argmax),
		.clk (clk),
		.rst (rstCosElement));
    end
endgenerate

reg [1 : 0] state;
always@(posedge clk)begin
	if (!rstCosElement)
		state <= INIT_ST;
	else begin
		case (state) // synopsys parallel_case
		INIT_ST:begin
					done <= 0;
					j <= 0;
					distance <= N;
					bestMatchID <= 0;
					if (argmax)
						state <= CNT_ST;
					else
						state <= INIT_ST;
				end
				 
		CNT_ST: begin
					if (distances[j] < distance) begin
						distance <= distances[j];
						bestMatchID <= j;
					end
					j <= j + 1;
					if (j > NUMLANG_MINES_1)
						state <= DON_ST;
					else
						state <= CNT_ST;
				end
				
		DON_ST: begin
					done <= 1;
					//if (argmax)
					//	state <= INIT_ST;
					//else
					state <= DON_ST;
				end

		endcase
	end
end

always @(posedge clk) begin
	if (!rst) begin
		langVectorsMem[ 0] <= textVector;
		langVectorsMem[ 1] <= textVector;
		langVectorsMem[ 2] <= textVector;
		langVectorsMem[ 3] <= textVector;
		langVectorsMem[ 4] <= textVector;
		langVectorsMem[ 5] <= textVector;
		langVectorsMem[ 6] <= textVector;
		langVectorsMem[ 7] <= textVector;
		langVectorsMem[ 8] <= textVector;
		langVectorsMem[ 9] <= textVector;

	end
	else begin
		langVectorsMem[ 0] <=10000'b0001000000100101000001101000111010100000000001011100100101110010110011011110011100000000000100000000100000101110101011101101000001110001010101111011110001100111011101011010010010010110100100100010000101111101010100100010001000101111001000100110001100000110000011011011110100111001011010000011101111010100000111100011111100001110010010011101011101011000011011000011111111101010001001111111001000110100010011110101000001001010100100111011110111101011011110101010110100110011000100111001101011111101110010010100101011000000001000010111100011110000111101110010111100111010101101000111101010110110010000001101010101010101010111111100011110100010100011010101101001010101110100101011011100011111011001001100111101011101011101111111001110110100000111101101100000101010100110000110101000111110100010101111000101000011101101100101101110100000100010011110101110110010100111001001011001000101110001100010000101101011000111101111001100111110010101101110111001100110000001100111001100010110111100101110110110111111011000101100101111001001010110101000010100000010110011101100111010110110111100101110110110011011010011010100010000100100010111101101100110101001011100011011110010000110011001111111100101101101101010001000001100010111000110010101110100101111110010001110011001001010111110110001101100111010110111110101110100000111011101111010101011101110010011001010110101010011000101100001100111011011010011011010001000111011110011001101011001110110101011101101011111111111000010111000100000011001011010001001110110000001001100101010101011101000000000111010011111101001100110101011001001011111100111100110100111100011011111000101111011110100101000001011111101010010010111011000001010001101001010111101001011001110110011100011010100101101001000111100011110100100010100010000011111100101101000000101011010111101011100001111110111011010001101000100101110010111101111100111101000100011100001100010000011100010001001011100010100110000010001010100011100000101100100100001011011110101100111111111010010001110111001111110011001101001100101101111110001011101000100111110010010001000011001010111011000011000110001001000110001010101001111011000010001110000011010011101111101101001111100010100010010100011000110011010001111011110101000101011110011011000110100101111011100010100000000011111101011001011010000100111001110101111110000100110110101001010001001101011001101101000000001010111101000000011110000001011001001010101100110010100101111111111010110000000010010011101011101100100110111011110110110011110111001100010010011101101010111110001000110100111001110110011001100111000111010011101100011100100000001100110000110110000111100000101101111000100110000101100110011111100100001101010011101111110111011110010100111001010110011100011001010111011010101011111110110010100101100001010111101000010101011001011101111111011001110100011101110110010000110001100111101011011001011010100011010100010000010010110101011111100110000010110011001000001010010111010101001111101000101101100100111111100011110111101001111001101110101100000011001010010010100110111011101110111111110100010001111011101001001001101000010011110111101000100111110011000000011100111101111001010111111000001011110101001101001000100001011110100110110011011100100000101001111100101101110100011011011010010111100000011000001101100100010101100010101110100110001001111110010100110100000100110001010101001100110011001101000011011001000111011000110010100000110001101110101000011000000010001011011011110001101001101111101000001100011100100010011100110000111011100101100100001101111011110110111010010110101101101011100011000011101100101100111001111001100010000111111100101111001000011100000110100011000100010000111010100000000101101001111110000001001111111000001110101111100110000110000111110001000010101001111001100001110110111010000101101001100011101001101100100111011000100110000110011110111101101011101000100011011010010101011010000100001010110010010100100000101111101010111110110110011101000010010011101100100111101011111111110011010000010010001001111110101001111010001000100110100011011010110000110110110110001001110001001111000111111010010000011100010001001011000101101001011110110111101100010111110110010001000111011001010011010001010000001011000011000100000000011010111101101100111011001011001110001010100111101110001110110000101101011010010111011101000011000010011011101010100010110100001101011001101111101001011111000000010111001010101101101101100000000100111110011011010010010111111111101001100110110111010100110000000011101101111110111100001110010111100100111000101101011000001110111001011001111000111100010101010110101110101011111110111110101110100000010010001011110100011100010001011111000011001000000111000001000001100111011110000111101011010000111011001100001011011000100001100000000011110100000000011010101000111111000110011111100000100101000111100001101000101111110011001101111110011011111111101111111111000011111100110110001001100100101000111100010100010010111010011100100110110101011000100111001111010010000000011110100100000011110011101101110111111010001101110111001101000001001110000110010101010000100110110101001101110101011101110001000100101111000110010011101111000101010110000110010000000111000001101010010000001111111100010101111001000100111110101101011010111000010110000101111111000101110011001110010111011010110000101100001100010101101110001100011100000010110101100001000101011110001011011010110111000100010010101011010101111000001111110010010010010010000111111101101000010100000101010011101001100101000010110010110111001001010010110101101011110001110011110001110110001010011011111010100000111111001100001101111010010110111000000010101001010010101110111101011001111011001101111011000101100010000111000111011000100011001011101010011111111100010111101010111010001110011100101001000011101011111110010111101100000011000100011101001001100001011101000101011000100110101110111011011110110001000111011111101101110110000010111001011011000100010010100011111010011110101001101010011111100011101010000111110001011100010001100000011111100000011101100001010000010110010111000111111011111110000100101011011100000011010011100110101111011000000111011001010011110010010111110110100110010000010100011110001111100001001010011100101000110110101111010110110100010111000101011100011001100011000100011110110101010001100010110101001101001111001000011000011000010011101101100111100110111000101111100111001010011001100001100001100010000011110011000111000000101110101011111001000101101111100111110100001111100100100000100011010010110100011001100010101110111011101110101101110000011010000101111001001010001110010101010111100100101101111100111101110010101100101011110110010000110010110001110001110011000100001101110111000000000100110010001000111111010010110010111101010000100100001001001000001100010111111100111001001010001100000111000010001001100010100100010011010111101000011010111000101001101011101101010101111111000001010011110010110001001011010001111011100011011011010110101010110001110111000001110111110001111100001111110111001111010100011100111010001111100000011001101110100110101000010011111001011001010110010010110111110010101011011110011011111110100111101100000111010011011001010001001100000010101001000110001011110001010111001000110001010111101010101101101101110111010101010010101010001011100010110111111010001011111000001001110110111100011010111000111110111100100110110010111111111001001001101011010111000011001001110100100011101011111101010100011100001111001011111010000110110110110011000110001100101010111111001110101101001110011001111110010101101110110000110110101011010011110000001010001110000010110100000100011110011100000000000110010111101110101001111100100011000110111100000100111000010000000001101111101001011001100011110100110111100010101111110000010011001010101100011011111110110010111011000001111101100100010101011100000111001001011101010000001000100001001101010101100101110100010100001011001001000001001001111111001100101001000111010100100001000110011010110100010010010000110101101100111001010110001010010011010110100010001011010011001110111111011110110000011101000110000010000000110010000011000000101111001010000011011111001100010000010011110101010000000011011100100110110111011011001011110100110010101101110011000010110011100110100000100111110110001101001011111101100110100101011010001011110000011000011010101011110000000100000000011000000011111010000110111010011100101010100111110010100000001000010001001110101010011010110010110001110101101110011010011101011000010010001100000110010011111001001100000111110011100110111000010011111111010110000000001000110110011000110001011011100001101001010011010000000001110111111110001111101001010001000100111111110001011110100111010001100011000011111101011100000100010010010010111010000100101110011000000011111110110111111111000101111010011010110101000011100111001001111110111001001101011010000101010001011001011101110010100100101101101110111110111110010100110101111010001110000000010011000100011111111111100001001011010110011101101101010110011101111111110100110110011000111001110000111010110010100011101100110011000011001000010011010011101010010100000001110111010000111110110011101010110001100010100010001100010100101000011001100011010001111100111000001100100010111111111010101110110000011010010101010100111010000000101000101010000111010011000001110110111111010111000001010000111111111001000111100011110000011000001001010110111101110101100000010110111010010001000111111101010111100010101110101011000000011001011101000110000010011000000111011100100111111101000100001010010100000111001000000111101100111010000111111011111110111100100001101000000011011010100110100111111010011010111110010100110110000000001011011111110011111011011011111110111011110001111101001011010001100110010001100110000110110001111010010010100100011011000110011100110110100000010000101001010111101111101010110100011100101000000110111000000001000101001100011110011100001110111001010110010101011100011011000011100111001001100111000001111100011000000110111011111011001001010000111100010110010111111110100011110011111000011111111011111111001101011011001; 
		langVectorsMem[ 1] <=10000'b0001000000100101010001101000111010100000000001011100110101110010110011011110011110000001000100000000100000101110101011101101000001110001010101111111110001100111001101011010010010010110100100100010000101111101010000100010001000101111001000100110001100000110000011011011110100111001011010000011101111010100000111100011011100111110010010011101011101011000011011000011111111101010001001111111001000110100010011110101000101001010100100111011110111101011011100101010110100110011000100111001101011111101110010010100101011000000001000010111100011010000111101110010111100111010111101000111101010110110010000001101010101010101010111111100011110100010100011010101101001010111110100101001011100011111011001001100111001011100011101111101001110100100000111101101100000101010100010000110101000111110100010101111000101000011001100100101101110000000100010011110101110110010110111001011011001000101110001100010000001101010000111111111001100111110010101101110111101100110000001110111001101010110111100101110110110111111011000101100101111001001010110101000010100000010110011101100111010110110111100101010100110011011010011010100010000100101010111101101100110101001011100011011110010000110011001111110100101101101101010001000001100010111000110010101110100101111110010001110011001001010111111110001101100111010110111110101110100000011011101111010101011101110010011001010111101010011000101100001100111011011010011011010001000111011110011001101001001110110101011101010011111111101000010111000100000011001011010001001110110000001001100101011101011101000000000111010011011101001100110101011101001011111100111100110100111111011011111000101111011110100101000001011111101010000010111011000001010001101001010111101001011001110110011100011010100101101001000111100011110100100010100011000011111100101101000000101011010111101011100010111110111011010001101000100101110010111100111100111101010100011100001100010000011100010001001011100010101110000010001010100111100000101100100100001011011110101100111111111010010001110111001111110011001111001100101101111110001011101000100111110010010001000001001010111011000011000110001001000110001010101001111011000010001100000011010011101111101101001111100010100010010100111000111111010001111011110101000101011110011011000110000101111011100011100000000111101001011001111010000110111001110101111111000100010110101001010001001101011001101101010000000010111101000000011110000001011001001010101100110010100101111111011010110000000010010011101001101100100110111011110110110011110111001100010010011101101010111110001000110100111001110110011001100111000101010111101100011100100000001100110000110111000111100000101101111000100110000101100110011111100100001101000011101011100111011100010100111001010110011100011001010111011010101011111110111010100101100001010111101000010101011001011101111111011011110100011101110110010000110000100111101011011001011010100011010100010000010010110101011101110110000010110011001000001010010111010101001111101000101001100100111111101111110111100001111001101110101100000010001000010000100110111011001110111111110100010001111011100001001001101100010011111111101000100011110011000000011100111101111001010111111000001011110101001101001000100001011110100110110011011100100000101001111100101101110100011111011010010111100000011000001101100100010101100010101110100110001001111110010100110100000100110001010101001100110011001101010011011001000111011000110011100000010001101110111000011000000010001011011011110001101001101111101000001100011100100010001100110000011011100101100100001101111011100110111010010110101101001011100011000010101100111100111001111001100000000111111100101111001000011100000110100011010101010000111010101000000101101001111100000001001111111000001110101111100110000110000110110001000110101001111101100001110110111010000101101001100011101001101100100111111000100110000110010110111101101001101000100011011010010001011010000100001010110010010100100000101111101010111110110110011101000010010011101100100111101011111111110011010000010010101001111110101001111010001000100110100011010010110000110110110110001001110001101111000011111110010000011100010001001011001101101001011110110111101100110111110110000001000111011001010011010011010000001011000011001000000000011010111101101100110011001010001110001010100111101110001110110000101101011010010111011101000011000010011011101010100010110100001101011001101111101001011111000000010111101000101101101101110000000100111110011011010010010111110111101001100110100111010101110000000011101111111110111100001110010111100100111000101101011000001110111001011001111000011100010101011110101110101011111110111110101110100000010010001011110100011100010001011111000011001000000111000001000001100111011110000111101011010000111011001110001010011000000001100000000011110100000000011010101000111111001110011111100000100101000111100001101000101111111011001101111110011011101111101011101111000011111100110110001001100100101000111100010100010010111010011100100010110100011000100110001111010110000000011110101100000011110011101101110111111010001101110111001101000001001110000010000101010000100110110101001111110101111101110001000100101111000110010011101111000101010110000110010000010111000001101010010000001111111100010101111001000000111110101101010010101001010110000101111111000101110010001110010111011010110000101100001100010101101110001100010000000010111101100101000101011110001011011010110111000101010010101011010101111100001111110010010010010110000111110101101000010100000101010011101001100101000010110011110111001001010010110101101011110011110011110001110110001010011011111010100000101111001000001101110010010110111000000010101001010010101110111101011001111011001101111011000101100010000111000111011000100011001011101010011111111100010111101010111010001110011100101001000011101011111110010111101100000011000100011101001001100001011101000101011000100110101110111011011110110001000111011111101101110110000010011001011011000100010010100011111010011110101001101010011111101011101010000111110001011101010001101000011111100000011101100001000000010110010111000111101011111110000100101011011100000011010011100110100111011010000111111001010011110010010111110110100110010000010100011110001111100001001010011100101000110110101111010110111100010111000101011100011001100011000100011110110101010001100010111101001100001111001000011000011000010011101101100011100110111000101111100111001010011001100001100001100010000011110011000111000000101110101011111001000101101111100111110000001111100000100000100011010010110000011001100010101110111011101110101101110000011010000101111001001010001110010101010111100100111101111100111111110010101100101011110110010000110010110001110001110011000100001101110111000000001100110010001000111111010010110010111000010000100100001001001001001100010111111100111001001010001100000111000010001001100010100100010011010111101000011010111000101001101011101101010101101111000001000011110010110001001001010001111011100011011011010110101010110001110111010011110111110001111100001111110111001011010100011100101010001111100000011001101110100110101000010011111001011001010110010010110111110010101011011110011011111110101111101100000111010011011001010001001101011010101001000110001011110001010111001000110001010111101010101001101001100111010101010010101010001011100010110111111010001011011000001001110110111110011010111000111110111100100010110010111111111001001001111011000111000011001001110100100011101011111101010100011100001111001011111010000110110110110011000110001100101010111111001110101101001110011001111110010101101110110000110110101011110011110000001010001110000010110100000000011110001100000000000110010111101110101001111100100011000110111100000100101000010000000001101111101001011001100011110100110111100110101111110000010011001010101100011011111110010010111011000001111101100100010101011110000111001001011101011000001000100001001101010101110101110100010110001011001001000000001001111111001100101001000111010100100001000110011010110100010010010000110101101100111001000110001010010011010110100010001011010001001110111111011110110000001101000110000010000000110010001011000000101111001010000011011111001100010000010011111101010000000011011101101110110111011011001011110100101010101101110011000010110011100110100000100111110110001101001001111101100110110101011011001011111000011100011010100011110000000100000000111000010011111010000110111010011100101010100111110010100000001000010001001110101010011010110010110001110101101110011010011101011000010011001000000110010011111000001100000111110011100110111000010011111111010110000000011000110110011000110001011011110001101001010011010000000001110111111110001111101001010001100100111101110001011110100111010000000011000011111101111100000100010010010010111010000100101010011000000011111110110011111111000101101010011010110001000011100101001001111110111001001101011010000101010001011001010101110010100100101101101110111110111110010100110101111010101110000000110011001100011111111111100001001011010110011101101101010110011101111111110100110110011000011001110000111010110010100011101100110011000011001000010011010011101010010100000001110111010000111110110011101010010001000010100010001100011100101000011001100011010001111100111000001100100010111111111010101110110000011010010101010100111010000000101000101010000111010011000001110110111111010111000001010000111111111001000110100011110000011000001001010110111101110101100000010110011010010001000111111101010111100010101110101011000000011001010101000110000010011000000111011100100111111101000100001010010100100111001000000111101100111010000111111011111110111100100001101000000011011010100110100111111011001010101110010100110110000000001011011111110011111011011011111110111011110001111101000011010001100110010001100110011110110001111010010010100100011011001110011100110110100010000000101001010111101111101010110100011100101000100110111000000001000101001100010110011100001110111001010111010101010100001011100011100111001001100111000001111100011000000110111011111011001001010000111100010110110111011110110011110011101100011111111011111111001101011011000; 
		langVectorsMem[ 2] <=10000'b0001000001100101010001101000111011100000000001011100100101110010110111011110011100000001000100000000100000101110101011101001000001110001010101111011110001110111001101011010010010010110100100100010000101011101010000100010001000101111001000100110001100000110000011011011110110111001011010000010101111000101000111100011111100011110010010011101011101011000011011000011111111101010101001111111001000110100010011110101010001001010100000111011110100101011011100101010100100110011000100111001101011111101111010010100101011000000001000010111100011010000111101110010111100111010101101000111101010110110010000001101010101010101010111111100111110100010100011010101101001010101110100101011011100010111011001001100111101011101011101111111001110100000000011101100100000101010100110000110101000111110110010101111000101000011101100100101001110100000100000011110001110110010100111001001011001000101110101100010000101101011000111111111001100111110010101101110111101110110000001110111001101010110111100100110110110111111011000101100101111001001010110111000010100000010110011101100111010110110111100101110010110011011010001010100010010100100010011101101100110101001011100011011110010100110011001110111100101101101101010001000001100010111000110010100110100111111110010001110011000001010111111110001101100011010110111110101110100000011011101111010101110101110010011001010111001010011000101100001100111011011010011011010011000111011110001001101011001110110101011101101011111111111000010111000100000011001011010001001110110000001001100101011101011101000000000111010001011101001100110101011111001011111100111100110100111111011011111000101111111110100101000001011111101000000010111011000001110001101001010111101001011001110110011100011010100101101001000111100011110100100010100011000011111100101101000000101011010111101011100010111110111010010001101000100101110010101101111100111101000101011100001100010000011100010001001011100010101110000010001010100011100000101100100100001011011110111100111111111010010001110111001111110011001101001100101101111110001011101100100111110010010001000001001010111011000011001110001001000110001010101001111011000010001100000011010011101111101101001111100010100010010101011000111011010001111011110101000101011110011011000100100101111011100011100000000011111101011001011010100100111001110101111010000100110110101011010001001101011001101101010000000010111101000000010110000000011001001010101100110010100101111111011010110000000010010011101011101100100110111011100110110011110111001100010010011101101010111110001000110100111001110110111001100110000101010111101100011100100000001100110001110110000111100000101101111000100110000101101010011111100100001101010011101011110111011100010100111000010110011100011001010111011110101011111110101010100101100001010111101000010000011001011101111101011001110100011101110110010000110001100111101011011001011010100011010100010000011010110101011111100110000010110011001000001010010111010101001111101000101011100100111111100011110111101001111001111110101100000011001000010010110110111011101110111111110110010001110011100001001001101100010011110111101001100011110010000000011110111101111011010111111000101011110101001101001000100001011110100110110011011100100000101001001100101101111100011111011010010111000000011000001101100100010101100010101110100110001001111110010100110100000100110001010101001000110011001001000011011001000111011000110011100000011001101110111000011000000010001011011011110001101001101111101000001100001100100010011100110000011111100101100100001101111010110110111010010110111101101011100011000010101100011100111001111001100010000111111100101111001000011100000110100011010100010000111010101000000001101001111110000001001111111000001110101111100110000110000111110001000010101001111101100001110110111010000100101001100011101001101100100111011010100110000110011110111101101011100000100011011010010001011010000100001010110010010100111000101111001011111110110110011101000010010011101100100111101011111111110011010000010010001001110110101001111010001000100010100011010010110000110110110110000001110001101111000111111110010000011100010001001011000101101001011110110111101100010111110110000001000111011001010011011011010000001011000011000100000000011010111101101100111011001010001110001010100111101110001010110000101101011110010111011101000011000010011011101010100010110110001101011001101111101001011101000000010111101010101101101101100000000100111110011011010010010111111111101001100110110111010100110010000011101100111110111000101110010111100100111000101101011000001110101001011001111000111100010101011110111110101010111110111110101110100000010010001011100100011100010001011111000010001000000111000001000001100111111110000111101011010000111011001110001010011000100001100000000011110100000000011010101001111111000110011111100000100101000111100000101000101111110011001101111110011011110111101111101111000011110110110110001001100100101000111100010100010010111010011100100110110100011000100111101111010010000000011111100100000011110011101101110111111010001100110111001101000001001110000010000101110000100100110101001101110101110101110001000100101111000110010011101111000101010110000110010000000111000001101010010000001111111100010101011101000000111110111100010010111001010110000101111111000101110011001110010101011010110000101100000000010101101110001100011100100010110111100101000101011110001011011010110111000101010010101010010101011000001111110010010010010010000110111101101000010100000101010011100001100101000010110010110111001000010010110101101011110011110011110001110110001011011011111010100000101111001100001101111010010110111000000010101001010110101110111101011001111011001101111011000101100010000111000111011000100011001011101010011111111100010111101010111010001110011100101001000011101001111110010111101100000111000101011101001011100001001101000101011000100110101110111011011110110001000011011111101101110110000010011001011011000100010010110011111010011110101001101010011111111011101010000111110001011100010001101000011111100000011101100001000001010100010111000111111011111110000100101011011100000011000011100110101111011000000111011001010011110010010111100110100110010000010100011110001111100001001010011100101000110110101111010110110100010111000101011100011101100011000100011110110101010001100010110101001101001111001000011000011000010011101101100111100110111000101111100111001010011001100001100001100010000011110011000111000000101100101011111001100101101111100111100100001111100100101000100011000010000100011001100010101110111011101110101101110000011011000101111001001010001110010101010111100101111101111100111101110010100100101011110110010000110010110001110001110011000100001101110111000000000100110000001000111111010010110010111000010000100100001001101100001100010111111100111001000010001100010111000010001001100010100100010011010111101000011010111000101001101011101101010101011111100001000011110010110011001011010001101111100011011011010110101010110001110111000001110111110011111100011111110111001111010100011100111010001111100000011000101110100110101000010011111001111001010111010010010111110010101011011110011011111110101111101100000111010011011001010001001100001010101001000110001011100001010111001000110001010111101110101001101101100011010101010010111010001011100010110111111010001011111000001001010110111110011010111000111110111100100100110010111111111001001001101011010111000011011000110100100011101011111101010100011100001111001011111010000110110110110011000110001100101010111111001100101101001110011001111110010101101110110000110110101011010011110000000010001110000010110100000100011110001100000000000110010110101110101001111100100011000110111100000100101000010000000001101111101001011001100011110100110111100110101111110000110111001010101100011011111110010010111001000001110101100100010101011110000111001001011101010000001000101001000101010101111101110110010110001011001001000000001001111101001100101011000101010100100001000110011010110000010010010000110101101100111001010110001010010011010110100110001011010011001110111111011110111000011101000110000010000001110010000010010000101111101010100011011111001100010000010011111101010000000011011100101110110111011011001011110100110010101101110011000010110011100110101000100111110110001101001001110101100110100101011010001011011000011010011010100011110000000100000000110000010011111000000110111010011000101010100111110010100000001000010001001110101010011010110010110001110101101110011010111101011000010010001000000110010011111001001101000111110011100110111000010011101011010110001000001000110110011001110011011011100001101001010011010110000001110111111110001111101101010001100100111111110001011110100111110000110011000011111100011100000100010010010010111010000100101010011000000011111110110111111111000101111010111010110101000011100111001001111111111001001101011010000101010001011011011101110010100100101101101110111110111110011100110101111010101110000000110011001100011111111111100101001011010110011101101101010110011101101111110100111110011001011001110000111010110010100011101100110011000011001000010011010011101010010100000000110111010000111110110011101010110001100010100010001100011100101000011001101011010101111100111000001100100010111111111010101110110000011010010101010100101011000000101000101010000111010011000001110110111111011111000001010000111111111001000110100011110000011000001001010110111101110101101000010110111010010001000111011101110111100010101110101011000000011001010101000110001010011000000111011100100111111101000100001010010100000111001000000111101100111010000111111011111110111100100001101000000011011010100110100111111010011010111110010100110110000000001011011111100011111011011011111110111011111001111101000011010001100111010001100110000110110001111010010010100100011011000110001100110110100000000000111001010111101111101010110100011100101000000110111000000001000001001100010110011100001110111001010111010100011100011011000011100111001001100111000001111100011100000110111011111011001001010000111100010110010111011110110011110011101100011111111011111111001101011011001; 
		langVectorsMem[ 3] <=10000'b0001000000100100010011101000111010100000000001011100110101110010110011011110011110000011000101000000100000101110101111101101000101110001010101111111110000100111001101011010010010010110100100100010000101011101010000100010001000101101001000100110001100000110000010011011110100111001011000000011101111011100000111110011011100111110010010011111001101011000011011000111111111101010001011111111001000111100010010110101000101001010101100101011110111101011011110101010111110110011000100111001101011111101111010010100101011000000001000010111100010010000111101110010111100111010111101000111101010110110010000001100010101010100010111111100011110100010100011010101101001010111110100101001011100011111111001001100111001011101011101111101001110000100000111101100100000101010100010000110101000111110101011101111000101000011001101100101101110000000100010011110100110100010110111000011011001000101110001100010000001101010001111101111001100111110110100101110111011110110000001110110001100010111111100100100110110111111011000101100101111001001010110110000010100000010110011101100111010110110111100101110100110011011010011110000010000100101010111101101100110101001011100011011110010000110011001111110100101101101101010101000001100110111000110010101110100111111110010001110001000001010111111110001101100111010110111110101100100100011011101111010101010101110010011001010111101010011000101100001100111011011000011011010101000111011110011001101101001110110101011001010011101111101000010111000101000011001011010001001110110000001001100101011101011101000100000111010011011101001100110101011111001011111100111100110100111111011011111000101111011110000101000001011111101010010010111011000001010001101001010111101001001001110110011100011010100101101001000111100011110000100010100011000011111100101101000000101011010111101011100011111110111110011001101000101101110010111100111100101101010100011100001100010000011100010001001001100010101110000010001010100111100000101100100100001011011110111100111111111010010001110111001111110011001111001100101101111110001011101000100111110010010011000011011010111011000011001111001001001010001010101001111011000010001100000011010011101111101101001111100010100010010100111000111111010001111011110101001101011110011011000100000101101011100011100000000111111001011001011010000110111001110111110011000100110110101001010011001101010001101101000000000010111101000000011111001101011001001010101100110010100111111111011010110010000010010011101011101100100111111010110110110011110111001100010000011101101010111110001000110100111001110110011001100111000101010111101100011100100000001100110001110111001111100000101101111001100110100101100110011111100100001100000011101011110111001100010100111001010110011100011001010101011010101011111110111010100101100001010111111000010101011001011101111101011011110100011101110110010000110000100111100011111001011010100011000100000001010010110101011101110110000010100011000000001010000111010101001111101000101101100100101111101111110111100001111101101110101100000010101000010000100110111011101110111111110100010001111011100001001001101100010011110101111000100011110011100000011100111101111000010111111000101011110101001101101000100001011110100010110011011100000000101001111100101101110100011111011010010111000100011000001101100100010101100010101110100110001001111110010100110100000100110001010101001100111010000001010011001011000111011000110011101000011001001110111000011000000010001011111011110001101001101111101010001100011100100010001100110000111011100001100100001101111001110110111010010110101101101011100011000010101100011100111001111001100000000111111100101111001000011100000110100011000001010000111010101000000101101001111100000001001111111000001010101111100010000110000111110000001110101001111001100001110100111010000101101001100011101001101100101111011000100110000110010110111101101001101000100011011010010001011010001100001010110010010100110000101111101010111110110110011101100010010011101100100111101011111111110011010010010010111001110110101001111010001010100110100011011010110100110110110100000001010001100111000011111010110000011000010101101011011101101001011110110111101100110111110110000001100111011001010011010010010000001011000011011100000000011010111101101100110011001000001111001010100111101110001110110000101001011010001111011101001011000110011011101010100010110100001101011001101111101001011111000000010111001000101101101101110000000100011110011011010010110111110101101001100110100011010101110000000010101111111110111000101110010111100100111000101101011000001110111001011001111001011100010101011110101110101010111111111110101110101100010010001011110100011100010001011111000010001000000111000001000001100111011110000111101011010000111011001100001011011000000001100000000011110100000000011010101000011111001110011111100000100101000111100001101000111111111011001101111110011011100111111111111111000011111100110110001001100000101000111100010100010010111010011100100010110100111000100110001111010110001000011111101100000011010011101101110111111010001101110111001101000001001110000010000101010000100100110101001111110101110101110001000100101111000110010011101111000101010110000110000100000111100001101010010000001011111100010101111001000010111110101101011010111000010110000101111111000101110010001110010101011010110000101100001000010101101110001100010000000000110111100101000100011110001011011010110111000101010010100011010101111100001111110010010010010110000111111101101000010100000101110011101001000101000010110011110111001001010010110101101011110011110011110001110110001010011111111010100000101111001000001100110010000110111000000011101001010010101110110101011001111011001101111111000101100010000111001111011001100011001011100010011111111100010111101010111010001110011100001001001011101011111110010101101100000011000101011101001001100001011111010101011000100110101110111011011110110001000011011111101101110110000010011001011011000100010010100011111010011110101001111010111111111011101110000111110001010100010001101000011111100000011101100001000000010100010111000111111011111110000100101011011100000011010011100110101110011010000111111011010011110010010111100110100110010000010100011110001111100001001010011100101010110110101111010110111100010111000101011100011001100011000110011110110101010001100010111101001100001101001000001000011000010011100101100011100110111000101111100111001010111001100000100001100010000011110011000111000000100100101011111001000101101111100111110000001111100000101000100011010010010100011001100010101100111011101110101101110000011010000101111001001010001110010101010111100100111101111100111111110010101100101111010110010000110010110001110001110011000100001101110111000000001100110010000100111111000010110010111000010000100100001001001001001100010111111100111001001010001100010111000010001001100010100100010001010111101000011010111000100001101111101101010101101111100001000011110010110011001001010001111011100011011011010111101010110101110111010011110110110001111100001111110111000111010100011100101010001111100010011001101111100110101000010011011001111001010110010010110111110010101011011100011011111110101111101100000111010011011001010001001101010010101101000110001011110000010111001100110001010101111010101101101001110111010101010010101010001011100010110011111010001011011000001001110110111110011010111000111110111100100010110010111101011001001000111011000111000111000001110100100011101011110101110100011110000111001011110010000110110110111011000110001100101010111111001110101101001110011001111110010101101110110000010110101011110011110001000010001010000010110100000000011110001100000000000110010111101110101001111100100011000010111100000100111000010000000001101111101001011001100011110100110111100110101111110000010011001010101100011011011110110010111011000001011101100100010101011110000111011001011101010000001000111001000101010101110101111100010110001011001001000000001001111011001100100011000101010101100001000110011010110100010010010000110101101100111001000110001010010011110110100010001011010001001110111111011110110000001101000110000010000000110010000011000000100111101010000011001111001100010000010011111101010000000111011100101110110111011011001011110100111010101101110001000010010011100110101000100111110110001101001001111101100110110111011011001011111000011100011010101011110000000100000000111000010011111000000110111010011100101010100111110010100000001000010001001110001010011010110010110001110101101110011010011101011100010011001100000110011011111001001101000111110011100110101000110011111111010110000000011000111110011010110011011011100001101001010001010000000001110111111110001111101001010001100100111111110001011110100111010010000011000011111111011100000100010010010010111010000100111110011000000111111110110111111111000111101010111010110001000011100101001001111110111001001101011010010101010001011001010101110010100100101101101110111110111110010100110100111010101110100010110011000100010111111111000001001011010110011101101101010110011101111111110100111110011000111001110000111000110010100010101100110011000011001001010011010011101010010100000000110111010001111110110111101010010001000010100010001100011100101000011001101011010001111100111000001101100010111111111010101110110100001010010101010100111010000000101000101010000111010011000001010110111111010111000001010000111111111001000111100011110000011000001001010010110101110101100000010110111010010001000110111101010111100010101010101011000001011001001101000110000010011000000111011100100111111101000100001010010100100111001000000111101100111000000111111011111111111100100001101000000011011010100110100011111011001001101110010100110110000000001011011111110011111011001011111110111011110001111100000011010001100110000001100110010110110001111010010010100100011011001100011100110110100010000000101001010111101101101010110100011000101000100110111000000001000001011100010010011100001110111001010111010100010100011011000011100111001001100111000001110100011000000110111011111011001001010000111100010110110111011110110011110011111000011111111011111111001101011011000; 
		langVectorsMem[ 4] <=10000'b0001000000100100000001101000111010100000000001011100100101110010110011011110001110000001000100000000100000101110101011101101000001110001010101111011110001100111001101011010010010010110100100100010001001111101010100100010001000101101001000100110001100000110000011011011110100111001011010000011101111010100000111100011111100101110010010011101011101011000011011000011111111101010101001110111001000111100010011110101000001001010101100111011110111101011011110101010100110110011000100111001101011111101111010010100101011000000001000010111100011110000111101110010111100111011101101000111101010110110010000001101010101010101010111111100011110100010100011000101101001010101110100101001011100011111011001001100111101011101011101111111001110100100000111101101100000101010100110000110101000111110110010101111000101010011101100100101101110100000100010111110100110110010100111000001011001000101110101100010000001101011000111111111001100111110110101101110111101100110100000110111001101010110111100101110110110111111011000101100101111000001010110101000010100000010111011101100111010110110111100101110100110011011010001010100010000100100010011101101100110101001011100011011110010000110011001110111100101101101101010101000001100010111000111010101110100101111110010001110001000001010111110110101101100101010110111110101110100010011011101111010101010101110010111001010111101010011000101100001100111011011000011011010001000111011110011001101011001110110101011001101011111111111000010111000100000011001011010001001110110000001001100101010101011101000000000111010011011101001100110101011111001011111100111100110100111100011011111000101111011110100101000001011111101010000010111011000001110001101001010101101001001001110110011100011010100101101001000111100011110100100010100010000011111100101101000000101011010111101011100001111110111011010001101000100101110011111101111100111101010100011101001100010000011100010001001011000010100110000010001010100011100000101100100100001011111110111100111111111010010001110111001111110011001111001100101101111110001011101000100111110010010001000001001010111011000011000100001001000110001010101001111011000010001100000011010011101111101101001111100010100010010100111000111011010001111001110101001101011110011001000110100101101011100010100000000111111101011001111010000110111001110101111110000100110110101011010001001101011001101101000000001010111101000000011110000101011001001010101100110010100101111111111010110000000011010011101001101100100111111011110110110011110111001100010010011101101010111110001000110100011001110110011001100111000101010111101100011100100000001100110000110110000111100000101101111000100010000101100110011111100100001101000011101111100111001110010100111001010110011100011001010111011010111011111110111010100101100001010111111000010101011001011101111111011001110100011101110110010000110001100111101011011001011010100011010100000000010010110100011101100110000010100011001000001010010111010101001111101000101001100100111111100011110111101001111001101110101100000011001000010000110110111011101110111111110100010001111011100001001101101100010001111111111000100111110011000000011100111101111001010111111000001011110101001101001000100001011110100110110011011100000000101001111100101101110100011111011010010111100000011000001101100100010101100010101110100110001001111110010100110100000100110001010101001100111011000101000011011001000111010010110011100000110001001110101000011000000010001011011011110001101001101111101000001100001100100010001100110000111011101101100100001101111011100110111010010110101101001011100011000010101100100100111001111001100010000111111100101111001000011100000110100011010100011000111010100000000101111001111110000001001111111000001110101111100110000110000111110001000010101001011101100001110100111010000101101001100011001001101100100111010010100110000110011110111101101001101000100011011010010001011010000100001010110010010100100000101111001011111110010110011101000010010001101000100111101011111111110011010100010010001001110110101001111010001010100110100011010010110000110110110110001001110001100111000111111110010000011100010001001011000101101001011110110111101100010101110110000001000111011001010011011011010000001011000001000100000000011010111101101100111011001001001111001010100111101110001010110000101001011010011111011101000011000010011111101010100010110100001101011001101111101001111111000000010111101010101111101101100000000100111110011011010010010111111111101001100110100111010100110010000011101101111110111100001110010111100100111100101101011000001110111001011001111000011100010101010110101110101010111110111110101110100000010010001011110100011100010001011111000010001000000111000001000001100111011110000111101011010000111011001110001011011000100001100000010011110100000000011010101000111111101110011111100000100101000111100001101000101111110011001101111110011011110111101011101111000011111100110110001001100100101000011100010100010010111010011100100010110101011000100111001111010010000000011110100100000011110011101101110111111010001101110111001101000001001110000110010101010000100100110101001111110101010101110001000100101111000110010011101111000101010110000110010000000110100001101010010000001111111100010101111001000000111110111101011010101000010110000101111111000101110011001110010101011010110000101100000100010101101110001100011100100010111101100001000101011110001011011010110111000100010010100011010101111100001111110010010010010010000111111101101000010100000101010011101001000101000010110010110011001001010010110101101011110001110011110001110110001010001011111010100000101111001000001101110110010110111000000011101001010010101110111101011001111111001101111101000101100010000111000110111000100011001011101010011111111100010111101010111010001110011100101001000011101011111110010111100100000111000100011101001011100001011101000100011000100110101100111011011110110001000111011111101101110110000010111001011011000100010011110011111010011110101001101010111111100011101010000111110001011100010001101000011111100000011101100001010001011110010111000111111011111110000100101011011100000011010011100110100111011000000111011001010011110010010111110110100110010000010100011110001111100001001010011100101000110110101111010110111100010111000101011100011001100011000100011110110100110001100010110101001101001101001000001000011000010011100101100111100110111000101111100111001010011001100000100001100010000011110011000111000000100110101011111001000101101111100111110100001111100100101000100011010010110100011001100010101110111011101110101101110000011010000101111001001010001110010101010111100100101101111100111101110010100100101011110110110000110010110001110001110011000100001101110111000000001100110000001000111111000010110010111100010000100100001001001000001100010111111100111001001010101100000111000010001001100010100100000011010111101000011010111000101001101011101101010101011101000001010011110110110001001011010001111011100011011011010110101010110001110111010001110111110001111100001111110111000111010100011100101010001111100000001001101110100110101000010011111001001001010111010010110111110010101011011110011011111110100111101100010111010011011001010001001110000010101101000110001011110001010111001100110001010111101110101001101101100011010101010010101010001011100010110111111010001001011000001001110110111110011010111000111110111100100010110010111111011001001001101011000111000011010001110100101011101011111101011000011100000111001011110010000100110110110011000110001100001010111111001110101101001110011001111110010101101110110000110110101011010011110000001010001010000010110100000100011110011100000000000110010111101110101001111100100011000110111100000100111000010000000001101111101001011001100011110100110111100010101111110000010011001010101100011011111110010010111011000000111101100100010101011100000111001001011101010000001000100001001101010101110101110100010100001011001001000001001001111111001100101001000101010100100001000110011010110100010010010000110101101100111001010110001010010011010110100010001011010011001110111101011110110000011101000110000010000001110010000011000000100111011110000011011111001100010000010011111101010000000111011100100110110111001011001011110100101110101101110011000010110011100110000000100111110010001101000011111101100110100101011011001010110000011010011010101011110000000100000000011000000011111010000111111010011100101010100111110010100000001000010001001110001010011010110010110001110101101110011010011101011000010011001100000010010011111001001000000111110011100110111000010011111111010110000000001000110110011001110011011011100001101001010011010000000001110111111111001111101001010001100100111101110001011110100111110000000011000011111101111100000100010010010010111010000100001110011000000011111111110111111111000101111010011010110101000011100101001001111110111001001101011000000101010001001001010101110010100100101101101110111110111110010100110101111010101110000000110011100101010111111111100001001011010110011101101101010110011101111111110100111110011000011001110000111010110010100011101100110011000011001000010011010011101010010100000001110111010000111110110011101010110001000010100010001100011100101000011001100011010001111100111000001100100010111111111010101110110000011010010101010100101011000000101000101010000111010011000001110110111111010111000001010000111111111001000110100011110000011000001001010110111101110101100000010110111010010001000111011101110111100010101110101011000000011001011101000110000010011000000111011100100111111101000100001010010100000111001000000111101100111010000111111011111110111100100001101000000011011010100110100111111010011010111110011100110110000000001011011111100011111011011011111110111001110001101100000011010001100110010001100110000110110001111010010010100100011011001110011100110110100000000000101001010111101101101010110100011100101000000110111000000001000101011100011010011100001110111001010111010101011100011011100011100111001001101111000001111100011000000110111011111011001001010000111100010110010111111110110011111011101101011111111011111111001101010011001; 
		langVectorsMem[ 5] <=10000'b0001000000100101000001101000111010100000000001011100110101110010110011011110011110000010000100000000100000101110101111101101000001110001010101111111110001100111011101001010010010010110100100100010000101111101010000100010001000101111001000100110001100000110000011011011110000111001011010000011101111011100000111100011011100101110010010011101011101011000011011000011111111101010001011110111001000111100010011110101010001001010101100111011110101101011011100101010110100110011000100111001101011111101110010010100101011000000011000010111100011010000011101110010011100111011111101000111101010110110010000001101010101010101010111111100111110100010100011010101101001010101110100101001011100011111011001001100111001011101011101111101001110000100000111101101100000101010100010000110101000111110100011101111000101000011001101100101101110100000100000011110101110110010110111011001011001000101110001100010000001101011000111101101001100111110011101101110111001110110000001110111001100010110111100101100110110111011011000101100101111001001010110111000010100000010110011101100111010110110111101101010010110011011010011010100010000100101010011101101100110101001011100011011110010000110011001111110100101101101101010101000001100010111000111010100110100101111110010001110011001001010111110110101101100111010110111110101110100000011011101111010101011101110010011001010111101010011000101100001100111011011010011011010101000111011110001001101101001110110101011101100011111111111000010111000101000011001011010001001110110000001001100101011101011101000100000111010001011101001100110101011011001011111100111100110100111111011011111000101111111110100101000101011101101010000010111011000001010001101001010111101001011001110110011100011010100100101001000111100011111100100010100010000011111100101101000000101011010111101011100011111110111010010001101000100101110010111101111100111101010100011100001100010000011100010001001001100010100110000010001010000011100000101100100100001011011110111100111111111010010001110111001111110011001111101100101101111110001011101000100111110010010001000011001010111011000011000110001001001110001010101001111011000010001100000011010011101111101101001110100010100011010100111000110111010001111011110101000101011110011011000100100101111011100010100000000011101001011001011010100100111001110101111111000100010110101001010011001101011001101101010100000010111101000000010111000000011001001010101100110010100101111111011010110000000010010011101011001100100110111011111110110011110111001101010010011101101010111110001000110100111001110110011001100111000101010111101100011100100000001100110001110111001111100000101101111000100010000101100110011111100100001100000011101011100111001100010100111000010110011100011001010111011010101011111110111010100101100001010111101000010101011001011101111111011011110100011101110110010000110000100111100011011001011010100011010100000000010010110101011101100110000010110001001000001010010111010101001111111000101001100100111111101111110111101001111001101110101100000010101010010010100110111011101110111111110100010001111011100001001001101100010010110111001000100011110011000000011100111101111000010111111000101011110101001101101000100001011110100110110011011100100000101001111100101101110100011111011010010111000010011000001101100100010101100010101110100110001001111110010100110100000100110001010101001100110011000001010011011001000111011000110011101000010001001110101000011000000010001011011011110001101001101111101000001100011100100010011100110000111111100101100100001101111011110110111010010110101101001011100011000011101100111100111001111001100000000111111100101111001000011100000110100011010101010000111010101000000100101001111110001001001111111000001010101111100110000110000110110001000010101001111101100001110100111010000100101001100011101001101100100111111000100110000110011110111101111001101000100011011010010101011010001100001010110010010100100000101111101010111110110110011101100010010011101000100111101010111111110011010010010010111001111110101001111010001010100110100011010110110000110110110110001001010001101111000011111010010000011100010001001011001101101001011110110111101100110111110110000001000111011001010011011011010000011011000011001100000000011010111101101100111011001010001110001010110111101110001010110000101101011110010111011101000011001010011111101010100010110100001101011001101111101001011111000000010111101000101101101101100000000100111110011011010010010111111111101001100111110111011100110010000011101111111110111000101110010111100100111000101101011000001110101001011001111000011100000101010110101110101010101110111110101110100000010010001011110100011100010001011111000010000000000111000001000001100111011110000111101011010000111011001110001011011000000001100000000011110000000000011010101001011111100110011111100000100101000111100000101000111111111011001101101110011011110111111011101111000011111100110110001001100100101000111100010100010010111010011100100110110101011000100110101111010110000000011111101100000011010011101101110011111010001101110110101101000001001110000110010101010000100110110101001101110101111001110001000100101101000110010011101111000100010110000110000000000111000001101010010000001011111100010101111001000100111110111100010010111001010100000101111111000101110010001110010101011010110000101100001000010101101110001100011100000011110111100101000100111110001011011010110111000101010010101011010101111000001111110010000010010110000111111101101000010100000101110011101001100101100010110011110111001001010010110101101011110011110011110001110110001010011011111010000000111111001100001101110010100110111000000010101001011110101110111101011001111011001101101001000101100010000111000111011000100011001011101010011111111100010111101010111010001110011100101001000011101001111110010101101100000111000100011101001001100001001111000101011000100110101110111011011110110001000011011111101101110110000010011001011011000100010010100011111010011111101001101010111111110011101010000110110001011101010001101000011111100000011101100001000000010110010111000111111011111110000100101011011100000011010011100110100110011000000011111011010011110010010111110110100110010001010100011110001111100001001010011100101010110110111111010110111100010111000101011100111001100011000100011110110101110001100010110101001100001111001000011000011000010011101101100011000110111000101111100111001010011001100000100001100010000011110011010111000000100110101011111001100101101111100111110100001111100000101000100011010010100000011001100010101100111011101110101101110000011011000001111001001010001110010101010111100100110101111100111111110010100100101011110110010000110010110001110001110011000100001101110111000000000100110010001100111111010010110010111000010000100100001001001001001100010111111100111001001010001100010111000010001001100010100100010011010111101010011010111000100001101011101101010101101111100001000011110010110011001011010001111011100011011011010110101010110001110111010011110111110011111100101111110111001111010100011100111010001111100000011001101111100110101000010011011001111001010110010010100111110010001011011110011011111110101111101100010111010011011001010001001101011010101001000110001011100001010111001100110001010111101010001101101001110111010101010000011010001011100010110111111010001011011000001001110110111110010010111000111110111000100100110010111101111001001000111011010111000011001000110100100011101011111101010100011100001111001011111010000110110110110011000110011100101010111111001100101101001110011001111110010101101110110000110110101011010011110000000010001110000011110100000000011110001100000000000110010110101110101001111100100010000110111100000100111000010001000001101111101001011001100011110100110111100010101111110000010011001010101100011011111110110010111011000000111101100100010101011110000111011001011101010000001010100001001101010101110101110100010100001011001001000001001001111111001100100001000111010100100001000110011010110100010010010000110101101100111001001110001010010011010110100010001011010011001110111111011110111000001101000110000010000000110010000011000000100111001010000011001111001100010000010011111101010000000111011101101110110111001011001011110100111110101101110001000010110011100110100000100111110110011101001011111101100110100101011011001011111000011000011010100011110000000100000000111000000011111000000110111010011100101010100111110010100000001000010001001110101010011010110010110001110101101110011010011101011000010011001100000110010011111000001100000111110011100110111000010011011111010110000000011000110110011001110011011011100001101001011011010000000001110111111111101111101101010001100100111111110001011110100011010000110011000011111110011100000100010000010010111010000100101110011000000011111110110011111111000101101010001010110001000011100111001001101110110001001101011010000101010001011001010101110010100100101111101110011110111110011100110101111010101110000000010011100101011111111111000001001011010110011101101101000110011101111111110100111110011000011001110000011010110010100011101100110010000011001000010011110011101010010100000000110111010000111110110011101010110001100010100010101100010100101000111001100011010101111100111000001100100010111111111010101110110000011010011101010100011010000000101000101010000111010011000001110110111111010111000001010000111111111001000111100011110000011000001001010010111101110101100000010110111010010001000111011101010110100010101110100011000001011001011101000110000010011000000111011100100111111101000100001010010101000111001000000111101100111010000111111011111110111100100001101000000011011010100110100111111010001010111110010100110110000000001011011111100011111011011011111110111011110001111101000011010001100110010001100110011110010001111010110010100100011011000110001100110110100010000000101001010111101111101010110100011100101000000110101000000001000101001100010110011100001110111001010100010001010100011011100011100111001001100111000001111100011000000110111011111011001001010000111100010110110111011110110011110011111100111111111011111111001101011011000; 
		langVectorsMem[ 6] <=10000'b0001000000100101000001101000111010100000000001011100110101110010111111011110011110000010000100000000100000101110101011101101000001110001010101111010110001110111011101001010010010010110100100100010000101011101010000100010001000101111001000100110001100000110000011011011110100111001011010000011101111001100000111100011111100100110010010011100011101011000011011010011111111101010001111111111001000111100010011110101010001001010100100111011110101101011011110101010110100110011000100111001101011111101110010010100101011000000001000010111100011110000111101110010011100111011111101000111101010110110010000001101010101010101010111111100111110100010100011010101101001010101110100101011011100011111011001001100111001011101011101111111101110100100000111101101100000101010100010000110101000111110100010101111000101010011011100100101101110000000100000011110101110110010110111001001011001000100110001100010000001101011000111101101001100111110011101101110111001100110000001110110001100010110111100100100110110111011011000101100101111001001010110110010010101000010110011101100111010110110111100101010010110011011010001010100010000100100010011101101100110101001011100011011110010100110011011111110100101101101101010101000001100010111000111010101110100101111110010001110011001001010111110110001101100111010110111110100110100000011011101111010101111101110010011001010111101010011000101100001100111010011010011011010101000111011110001001101111001110110101011101101011111111111000010111000100000011001011010001001110110000001001100101011101011101000000000111010001111101001100110101011011001011111100111100110100111111011011111000101111111110100101000001011111101000000010111011000001010001101001010111101001011101110110011100011010100100101001000111100011111100100010100010000011111100101101000000101011010111101011100011111010111010010001101000101101110010111101111101111101000100011100000100010000011100010001001001100010100110000010001010000011100000101100100100001011011110111100111111111010010001110111001111110011001101101100101101111110001011101000100111110010010001000001001010111011000011001110001001000110001010101001111011000010001100000011010011101101101101001111100010100010010100111000110111010000111011110101000101011110011011000100100101111011100010100000000011111101011001011010000100111001110101111111000100110110101011010011001101011001101101000100000010111101000000011110000001011001001000101100110010100101111111011010110000000010010011101011001100100110111011101110110011110111001100010010011101101010111110001000110100111001110110011001100111000101010011101100011100100000001100110001110111001111100000101101111000100010000101111110011111100100001101000011101011110111011100010100111000010110011100011001010111011010101011111110111010100101100001010111101000010001011001011101111111011011110100011101110110010000110001100111100011011001011010100011010100000000010010110101011111100110000010110011001000001010010111010101001111101000101001100100111111100111010111101001111001101110101100000010101010010010100110111011101110111111110110010001111011100001001001101100010010110111001000101111110010000000011110111101111001010111111000001011110101001101101000100001011110100110110011011100100010101001111100101101110100011111001010010111000010011000001101100100010101110010101110100110001001111110010100110100000100110001010101001100110011000101000011011001000111011000110011101000010001001110101000011000000010001011011011110001101001101111101000001100011100100010011100110000111111100101100100001101111011110110111010010110101101101011100011000010101100011100111001111001100010000111111100101111000000011100000110100011010101010000111010100000000101111001111110001001001111111000001110101111100110000110000111110001001010101001111101100001110110111010000100101001100011101001101100100111111100100110000110011110111101111001101000100011011010010101011010001100001010110010010100110000101111101010111110110110011101000010010011101000100111101011111111110011010010010010111001111110101001111010001000110110100011010110010000110110110110001001110001001111000111111010010000011100010001001011001101101001011110110111101100110111110110000001000111011001010011011011010001011011000011001100000000011010111101101100111011001010001111001010100111101110001010110000101101001010010111011101000011000010011111101010100010110100001101011001101111101001011111000000010111001000101101101101100000000100111110011011010010010111111111101001100110110111011100110010000011101111111110111000001110010111100100111000101101011000001110101001011001111000011100010101010110101110101010101110111110101110100000010010001011100100011100010001011111000010000100000111000001000001100111111110000111101011010000011011001110001011011000100001100000000011110000000000011010101001011111100110011111100000100101000111100000101000101111111011001101111110011011110111101011101111000011111110110110001001100100101000111100010100010010111010001100100110110101010000100110101111010110000000011111101100000011110011101101110011111010001101110111101101000001001110000110010101010000100110110101001101110101111001110001000100101101000110010011101111000101010110000110000000000111000001101010010000001111111100010101111101000100111110111100010010111001010110000101111111000101110010001110010101011010110000101100001000010101101110001100011100100010110101100101000100111110001001011010110111000101010010101011010101111000001111110010000010010010000110111101101000010100000101110011101001100101100010110011110111001001011010110101101011110011110011110001110100001011011011111010100000101111001000001101111010100010111000000010101001011110101110111101011001111011001101111001000101100010000111000111011000100011001011100010011111111100010111101010111010001110011100101001000011101001111110010101101100000111000101011101001001100001011111000101011000100110101110111011011110110001000111011111101101110110000010111001011011000100010010100011111010011111101001101010011111100011101010000110110001011101010001100000011111100000011101100001000001010110010111000111111011111110000100101011011100000011010011100110100111011000000111111011010011110010010111110110100110010000010100011110001111100001001010011100101010110110111111010110111100010111000101111100111001100011000110011110110101110001100010110101001101001111001000001000011000010011101101100011110100111000101111100111001010011001100001101001100010000011110011010111000000100110101011111001100101101111100111110100001111100000100000100011010010110000011001100010101100111011101110101101110000011011000101111001001010001110010101010110100100100101111100111101110010100100101011110110010000110010110001110001110011000100001101110111000000000100110000001100111111010010110010111000010000100100001001001100001100010111111100111001001010001100010111000010001001100010100100010011010111100010011010111000100001101011101101010101111111100001000011110010110001001011010001101111100011011011010110101010110001110111010011110111110011111100111111110111001111010100011100111010001111100000011001101110100110101000010011011001101001010110010010110111111010001011011110011011111110101111101100000111010011011001010001001101001010101001000110001011110001010111001100110001010111101010101101101001100011010101010010111010000011100010110111111010000011011000001001110110111000010010111000111110111000100100110010111101111001001000101011010011000011001000110100100011101011111101110100011100001111001011111010000110110110110011000110001100101010111111001110101101001110011001111110010101101110110000110110101011010011110000000010001110000010110100000100011110001100000000000110010110101110101001111100100011000010111100000100111000010001000001101111101001011001100011110100100111100010101111110000010011001010101100011011111110110010111011000000111101100100010101011110000111011001011101010000001001100001001101010101110101110100010100001011001001000000001001111101001100101001000111010100100001000110011010110000010010010000110101101100111001001110001010010011010110100010001011010011001110111111011110011000001101000110000010000000110010000011000000100111001010000011001111001100010000010011111101010000000111011100101110110111011011001011110100111110101101110001000010110011100110100000100111110110011101001011111101100110100101011010001011111000011000011010100011110010000100000000111000000011111000000110111010011100101010100111110010100000001000010001001110101010011010110010110001110101101110011010011101011000010011001000000110010011111000001100000111110011100110111000010011011111010110000000011000110110011001110011011011100001101001011001010010000001110111111111001111101000010001100100111111110001011110100111010000110011000011111111011100000100010010010010111010000100101110011000000011111110010011111111000101100010001010110001000011100111001001111111111101001101011010000101010001011001010101110010100100101101101110111110111110010100110101111010101110000000010011001101011111111111000001001011010110011101100101000110011101111111110100110110011001111001110000011010110010100011101100110011000011001001010011110011101010000100000000110111010000111110110001101010110001100010100010101100010100101000011001100011010101111100111000001100100010111111111010101110110000011010011101010100001010000000101000101010000111010011000001110110111111010111000001010000111111111001000111100011110000011000001001010010111101110101100000010110111010010001000111011101010110100010101110100011000001011001010101000110000010011000000111011100100111111101000100001010010101000111001000000111101100111010000111111011111111111100100001101000000011011010100111100111101010001010111110010100110110000000001011011111110011111011011011111110111011110001101101001011010001100110010001100110011110010001111010011010100100011011000110001100110110100000000000101001010111001111101010110100011100101000000110111000000001000101001100010110011100001110111001010100010001010100011011100011100111001001101111000001111100011000000111111011111011001001010000111100010110110111011110110011110011111100111111111011111111001101011011000; 
		langVectorsMem[ 7] <=10000'b0001000001100101000001101100111010100000000001011100100101110010111011011110001110000010000000100000100000101110101011101101000101110001010101111011110001110111001101001010000010010110100100100010101101011101010100100010001000101111001000100110001100100111000011001011110000110101011010000011101111010100000111100011111100100110010010011100011111011000011011010011111111101010001011110111001000111100010011110101010001011010100100111011110110101011011101101010111100110011100100111001101011111101110010110100101011000000011000010111100011110000111101110010111100111010111101000111101010110110010100001101010101010101110111111100111110100010000011011101101101010111110100101001011100011111011001001100111001011101011101111101001110000000000011001101100000101010100010000110101000111110101010101111000101010011001101100101101110100000100010011110001110110010110111011011011001000100110101100010000101101011000111111101001100111110011100101110111001000110100001110110001100010110111101100110110110111011011000101100101111001001010000101000010100000010110011101000111010110110111100101110000110011011010011010100010000100100010011101101100110100001001100011011110010100110011011111110000101101101101010101000001100010111000111010100110100101111110010000110011000001010111110110001101000111010110111110011100100100111011101111010101101101110010011001010111101010011000101100001100111010011010011011010001000111011110011001101111001110110101011101000011111111101000010111000101000011001011010001001110110000001001100101110101011101000100000111110001111101001100110101011001001011111100111100110100111111011011111000101111011110101101000001011001101000010010111011000001110001101001010101101001011101110100011100111010100101101000000011100011111000100010101010000011111100101101000000101011010110101011100011111111111010011001101000101101110010111101011101110101010100011100000100010000011100010011001001100010100110000010001010000011100000101100101100001011011010011000111111111010010001110111001111110011011101101100111101111110001011101100100111110010010001000011001010111011000011000101001001000110001010101001111011000010001100000011010011101101101101001111100010100001010100111010110111010000111011110101000101011110011001000110000100111011100010100000000001111101011001011010100100111001110101111111100100110110100101010011011101011001101101010101000010111101000000011110000000011001001000101110110010101111111111011111110000000010000011101011001100100110111011101110110011110111001100010010011101101010111110001000110101111001110110011001100011000101010111101100011100100000001100110001110111001111100000101101111000100010000001111111011111100100001101000011101011100111111100010100111000010110011100011001010101011110101011111110100010100101100001010111101001010000011001011101111111001011110100011101110110010000110000100111100011011001111010100011010100010100011010110100011111100111000010110001001000001010010111111101001111101000101001100100101111111111110111101001111001101110101100000010101000010000110110111011101110111111110110010001111011100000000101101100011010110101001000100011110011100000011110111100111011010111111000101111110101001101001000100001010110100110110011111100000010101011111100101101111100011111011010010011000110011000001101000100010100100010101110100010011011111110010100110100000100100001110101001100110011001001000011011011000111011000111001100000100001001110101000011000000010001011111011111001101001101111101000001100011100100010011100110000011111001101100101001101111011100110111010010110101101101011000011000011101100001100111001111001100010000011111100101111000000011100000110100011010101010000111010101000000101111001111110000101001111111000001110101111100110010110000111110001001010101001011001100011111110111010000100101001100011101001101100100111110010100110000110010110111101111001101000100011010010010101011010001100001010110010010100110000111111101000111110010110000101000010010011001000100111101010111111110011110010010010111001111110101001111010001000110010100001010010110000110110110110001001110001001111000111111110010000011100010001001011000101101100011110100111101100110101110110000001101111011001010011011011010000010111000011001100000000011010111101101100111011001001001110001010100111101110001010110000101100011110010111011101000011001110011111101000100010110100001101011001101111101001011111000000010111101000101101111101100000000100111110011011010010010111110111101001100100010111011101110010000011101011111110111101101110010110100100111100101101011000001110111001011001111000111110000101010110101010101011101110111110101110100000000010001011110100011100010001011111000010000100000011000001000001100111011100000111101011110000011011111110001011011000100001000000000011110100000000011010101001011111100110011111100000100101000111100000101000100111111011001101101111011011110111111001101011100011110100110110001001100100101100101100010100010010111010001101100110110100011000100100001111010110000000011110100100000011010011101101110011111010001001110111001101000001001110000010010101010000100110110101011101110101011101110001100100101101000010010011101111000100010111000110010000101111000001101010010000001111111100010101111001000000111110111000010010111001010110000101111111000101110010000110010101011010110000101100001100010101101110001100011100000011111101100001000100111110001011011010110111100100010010101011010111111000001111110010000010010010000110111101101000010100010101010011101001100101100010110011110111000001010010110101101011110011110011100001110110001010011011111010100000111111001000001001111010100000111000000010101001011110101110111101011001110011101101101001000101100010000111000111011000100011001011100010011111111100010111101010111010001110011100101011000011101011111110010101101100000111000101011101001001100001011111010101011000100110101110111011011110100001000101011111101101110010000010011000011011000100010010100010111010011110101001101010110111110011101010000110110001011101010001101110011111100000011101100001000000011100010111000111111011111110000100101011011100000011011011100110100111011000000111011001010011110010010111110110100110010000010100011110001111100001001010011100101010110110111111010110111100010111000101111100111101100011000100011110110101110001100010110111000101001111001000011000011000000011101101100011000100111000101111100111001010011001100000101101100010000011110011010111000000101110101111111001100101101111100111110000001111101000101001000011000010100000011001100010101110111011101110101101110000111011000001011001001010001110010101010111100101110101111100111111110010100100101010110110010000110010110001110001110011000100001101110101000000001100110000001100111111010010110010101000010000100110001001101001001100010011111100111001001010001100010111000010001001100010100100010011010111101010011010111000100001101011101101010101011001100001000011110010110011001011010001111011000011011011000100101010110101110111010011110111110011111100111111110111001111010110011100111010001111100000011001101110100110101000010011001001001001010110010010110111111110001011111100011011101110101111101100010111010011011101010001001101011010101001000110001011100000010111001100110001010111101110101001101001100011010101010001111010001011100010110111111010001001011000001001010110101100010010111000111110111001110100100010111101110001001001101011001111000011011000110100110011101011111101111100011110001111010011111010000100110110110011000110001100001010111111001110101101001100011001111110010101101110110000110110101011010011110000000010001110001011110100000100011110011100000000000110010110111110101001111100100011000010111100000100111000010001000001101111101001011001100011110100110111100010101111110000110011011010101100011011111110110010111011000001110101100101010101011110010111011001011101000000001001110001001101010101110101110100010100001011001001000000001001111111001100100001000001010100100001000110011010110000010110010000110101101100111001010110001010010011010110100010001011010011001110111111011110010000001101000110000110000000110110010011000000100111101010000011001111001101000000010011111101010000000011011100100110110111011011011011110100111110101101110001000010110011100110100000100111110110011101001001111101100110110101011010001011111000011000011010100011110010000100000000111000000011111000000110111011011100101010100111110010100000001010010001101110101010011010110110110001110101101110011010011101011000010011001100000110010011111000001100000111010011100110111000010011001111010110001100011000110110011001110011011011100001101001011001010010000001110111111111101111100000010001100100111111110001011110100011010000110011000011110110011100000100010000010010101010000100101110011010000011111111010011111111000111111010001010110101000011100101001000111111011101001101011000000101011001001001010101110010100100101101101110011110111110011100110101111110101100010000010011100101011111111111000000001011010110011101100101000110011101111011110100110110011001111001110000011110110010110011101100110011000001001000010011110011101010010100000000110111010000111110110001101010110001100010100010000100010100101000011101100011010101101100111000001101100010111111111000101110110000011010010101010110011010001000101000101010000011000011000101110110111111011111000001011000111111111001000111100011110000011010001001010010111101110101100100010111111010010001000111011101010110101010101010100011001001010001011101000100011010011000000111011100100111101111000000001010010101000111001000000111101100111000000111111011111110111100100001101010000011011010100111100110111010011010101110010100110100000000001011011111100011111011011011111110111011110001101100001011010001100111010001101110011110010001111010011010100100011001000100001100110110100010000000101001010111001111101010110110011100001000100110111000000001000101001100011110011100011110011001010100010001010100011011100011100111001001101111000001111100011000000111111010001011001001010000111100010110110111011110100001110010111000011111111011111111001101011011011; 
		langVectorsMem[ 8] <=10000'b0001000001100101000001101000111011100100000101011100110101110010111110001110001110000001000100000000100000111110101111101001000001110001000101111011110001100111011101011010010010010110100100100010000101111101010100100010001000101101001000100110000110000110000011001011110110110001011010000011101111000101000111100011011100001110010010011101011101011000011011010011111111101010101001011111001000111100010011110101000001011010100100111011010111101011010110101010100110110011100100111001101011111101110010011100101011000000001000010111100010110000111101110010111100111011101101000111101010110110010000001101010101010101010111111100011110100010100011000101101001010101110100101011011100011111111001001100111101011100011101111111001110110100000011101111100000101010100110000110101000111110110010101111000100010011001100100101101110100000100010011110101010110010110111001001011001000101110001110010000101101011000111111111001100111100010101100110111101100110000000100111001101010111111100111110110110111111011000101100101111000001010110100010010100000010100011101100111010110110111100101110110110011011010011010100110000100100010111101111100110101001011100011011110010100110011011110111000101101101101010001000001100010111000110010101110100101111110000001110001000101010111110110101101100111010110111110001110100010011011100111010101010101110010011001010110101010011000101100001100111011011010111011010001000111011110011001101011001111110101011101111010001111111000010111000100000011001011010001001110110000001001100101010001011101000000000111010011111101011100110101011001001010111100111100110100111010011011111100101111011110100111000001011011101010010010111010000001010001101001010111101001011001010110011000011010000101101001000011100011110100100010100010000011111000101101000000101011010011101011100001111110111011010011101000100100110011111101111100111101100100011101001100010000011100010001001001100111100110000010001010100011100000101100100100001011011110111100111111111010010001110111001111110011001101001100101101111110001011101000100111110010010001000001001010101011000011000110001001000110001010101001111011000010011110000011010011101111101101001111100010100011010001011000110011010001101011110101000101001110011001000110000101101011100010100000000111101101011000011010000110111001110111111110000100110110101001010001001101011001101101000100000010111101000000011110000100011001001000101100110010100101111111011010110000000011010011101011101100100111111011110110110111110111001101010000011101101010111110001000110000111001110110111001100110000101010011101110011100100000001100110000110110000111100000101101111000100110000101100110011111100100001101000001101111110111011110011100111001010110011100011001010111011110101011111110110010100101110001010111111000010101011101011101111111011001110100011101110110010000110001100111101011111001111010100011000100010001110010110101011111110110000010100011000000001010010111010101001111101000101001100100111111100011010111101001111001101110101100000011001010000000110110111011101110111111110100010001111011101001001001101100011001111111101000100111110011001000011101110001111001010111111000001011110101001101001000100001011110100110010011011100000000101001011100101101110100011111011010010111100000010000001101100100010101100010101110100110001001111110110100110100000100110001010101000100110011001001000011011001000111011000110010110000110001101110101000011000000010001011011011110101101001101111101000001100001100100010011100110000011111100101100100011101011011100110111000010110101101101011100011000010101100001100111001111001100010000101111100001111001000011100000110100011010000010000111010100000000101101001111110000001000111111000001110101111000110000110000101110001001010101001011101100001110100111110000101100001100001101001101100101111111000100110000110011110111101001011100000100001011010010101011010000000001010110010010100110000101111001011111110110010001101000010010011001000100111100010111111110011010100000010100001110110101001111010001010110010100011011010110000110110110110000001110001000111000111111110010000011100010001001011001101101001011110110111101100010111110110010001001111011001010011011011010000001011000001000000000000011010111101101100111011001011001110001010100111101100001110110000101101011010010111011101000011000010011011101010000010110100001101011001101111101001011111000010000111001000101111101101100000000100101110011011010010010111111111101001100110100011010110110010000011101101111110111100001110010110100100111100101101011000001110111001011001011000111100000101010110101110101011111110111110101110100100010010001011110000011100010001011111000011001000000110000001000001101111011110000111001011010000111011111100001011011000000001100000000011110000000000011010101000111111001110011111100100100101000111100001101000101110111011001100111110011011111111101011111111000011111100110110001001100000101000011100011100010010111010011100110110110101011000100110001110010010001000011110100100000011110011101101111111101010011101110111001101000001001110000110000101010000000100110101011111110101111001110001000100101111000111010011101111000101010110000110010000010111100001101010010000001111111100010101111001000100111110111101010010111001010110000000111111000101110011001110010111011010110000101100001100010101101110001100011100000010111101100001000101011110001011011010100111000110010010101011010101111100001111110010100010010010000111111101101000010100010101010011101001100101000010110110110111001001010010110101101010010001110011100001110010001010001011111010100000101111001000001101111110010110111000000010101001010110101110111101011001111011001101111001000101100010000111000111111000100011001011101010011111111100010111101110111010001110011100101111000111101011111110010111100100000111000101011101001011100001011101000101011000100110101110101011011110110001000101011111101101110110000010111001011011000100010110100011111010011110101001111010011111100011111110000111110001011100010001100000011111100000011101100001010000010110010111000111101011111110000100101011011100000011010011100110101111011000000111011001010011110010010111110110100010010000010100011110001011100001001010011100101000110110101111010110110100010111000101111100011001100011000110011110110100010001100010110101001100001111001000011000011000010011101101100010100110111000101111100111001010011001100001100001100010000011110011000111000000101110101011111001100101101111100111111100001111100001100000100011010010110100011001100010101110111011101110101101110000011011000101111001001010001110010101010110100100111101111100111101110010101100101011110110010000110010110001110001110011001100001101110111000000001100110010000001111111110010110010111101010000100100001001001000001100010111111100111001000010001100000111000010001001100011100100010011010101101000011010111000101001101011101101010101011101000001110011110010110001001011010001101011100011011011010110101010110001110111001001110110110001111100011101110111000011010110011100110010001111100000011001101110100110101000100011111001001001010110010010010111111010101011011110011001111110100111101100000011010011011001010001001100010010101101000110001011110001010111001000110001010111101110101001101101100111010101010010001010001011100010110111111010001001111000001001110110110100011010111000111110111000100010110010011111010001001001101011010111000011010001110100001111101011111111010100011100101111001011111010000110110110110011000110001100101010111111001100101101001110001001111110010101101110110000110110101011110011110001001010001010000010110000000100011110011100001000000110010110101110101001101100100011000110111100000100110000010000000001101111101001011001100011110100100111100010101111110000010011001110101100011011111110010010111011000000110101100100010101010100000111001001011101000000001001110001001101001101100101110100010100001011001001000001001001111111001100101011000011010100100001000110011100110000011010010010110101101100111001010110001010010011010110100110001011010011001110111101011100111000011001000110000010000000110010001011000000101111001010100011011111001100010000010011101101010000000011001101100110110111011011001011110100100010101101110011000010100011100110100000100111110110011101001011111101100110100101011010001010110000011110011010101011110000000100000000011010000011111010000110111011011100101010100111110010100000001010010001001110101010011010110010110001110101101110011010111111011000010011000100000010011011111000001000000111110011100110111000010011111011010110000000111000110110011001110001011011110001101001010011010110000001110111111110001111101001010001000100111111010001011110100111110000010011000011111101111100000100010011010010111010000101111110011000000011111110110111111111100100111010011010110001000111100111001001111110111001000101011000000101010001001001010101110010100100101101101110111110111110010100110101111010101110010000110111000100010111111111100001001011010110011101101101110110011101101111110100110110011000111001110000111010110000100011101100110011000011001000010011010011101010010100000001110111010000111110110011101010010001000010101010000100010100101000010001100011110101111100111000001100101010111111111010101110110000011010011101010110101011000000101000101010000111010011000001110110111111010111000001010000111111111001000110100011110000011000001001010110110100110101100000010110011010010001000101111101010111100010101110101011000000011001010101000100000010011000000110011100100111111101000100001010010101000111001000100111101100111000000111111011111110111100100001101000000111011010100110100111111011011011110110111100110110000000001011011111110011111011011001101110111001110001111100001011010001100110010001101110000110110001111010110010100100011011001110001100100110100000000000101001010111001111101010110100011100001000000110111000000001000101001100011111011100001110111001010110010101011110001011000011100111001001100101000001101100011000000110111011111011001001010000111100010110010111111110100011110010101000011111111011111111000101001011001; 
		langVectorsMem[ 9] <=10000'b0001000000000101000001101000111011100100000001011100110101110010111111001110001110000001000100000000100000101110101011101001000001110001010101111011110001100111001101011010010010010110100100100010000101011101010100100010001000101101001000100110001100000110000011011011110100111001011010000011101111001101000111100011111100000110010010011101011101011000011011010011111111101110101001111111001000110110010011110101000001001010100100111011110111101011011000101010100110110011100100111001101011111101110010011100101011000000001000010111100011110000011101110010111100111011101101000111101010010110010000001101010101010101010111111100011110100010100011000101101001010101110100101011011100011111011001001100111101011101011101111111001110100100000111101101100000101010100110000110101000111110100010101111000101010010001100100101101110100000100010011110101110110010110111001001011001000101110001110010000101101011000111111111001100111110011101100110111001100110000000100110001101010110111100101110110110111111011000101100101111101001010110101010010100000010100011101100111010110110111100101010110110010011010001010100110000100100010111101101100110101001011100011011110010000110011001110111000101101101101010001000001100010111000110010101110100101111111000000110011001001010111111110101101100111010110111110001110100000011011101111010101010101110010011001010111001010011000101100001100111011001000011011010001000111011110011001101011001110110101011101101011111111111000010111000100000011001011010001001110110000001001100101010101011101000000000111010011111101001100110101011001001011111100111100110100111011011011111000101111011110100101000001011001101010000010111011000001110001101001010111101001011001110110011000011010100101101011000111100011110100100010100010000011111000101101000000101011010111101011100011111110111011010001101000100100110011111101111101111101010100011101001100010000011100010001001011100010100110000010001010100111100000101100100100001011011110101100111111111010010001110111001110110011001101001100101101111110001011101000100111110011010001000001001010101011000011000110001001000110001010101001111011000010001110000011010011001111101101001111100010100010010000011000110011010001111011110101000101011110011001000100100101111011100010100000000011101101011001011010000110111001110111111110000100110110101001010001001101011001101101010000001010111101000000011110000001011001001000101100110010100101111111011010110000000010010011101001101100100111111011110110110111110111001101010000011101101010111110001000110100111001110110011001110111000111010011101100011100100000001100110000110110000111100000101101111000100110000101100110011111100100001101000011101111110111011100011100111001010110011100011001010111011110101011111110110010100101100001010111111000010101011001011101111111011001110100011101110110010000110001100111101011011001111010100011010100010100010010110100011101100110000010100011001000001010010111010101001111101000101001101100111111100011110111101001111001101110101100000011001010000000100110111011101110111111110100010001111011101001001101101100010011111111101001100111110010000000011100111001111001010111111000001011110101001101001000100001011110100110110011011100000000101001011100101101110100011111011010010111100100011000001101000100010101100010101110100110001001111110010100110100000100110001010101001100110011001101010011011001000111011000110010100000110001101110101000011000000010001011011011110001101001101111101000001100011100100010001100110000011111100101100100011101111011100110111010010110101101101011100011000011101100000100111001111001100010000111111100001111001000011100000110100011010100010000111010101000000101101001111110000001001111111000001110101111000110000110000111110001001110101001011101100001110100111010000101100001100011001001101100100111111000100110000110011110111101101011101000100001011010010101011010000100001010110010010100110000101111001011111110110110001101000010010011001000100111100010111111110001010100010010000001111110101001111010001010110110100011011010110000110110110110001001110001000111000111111110010000010100010001001011001101101001011110110111101100010101110110000001000111011001010011010011010000001011000011000000000000011010111101101100110001001010001111001010100111101110001110110000101101011010010111011101000011000010011111101010100010110100001101011001101111101001011111000000000111001000101111101101110000000100111110011011010010010111111101101001100110100110010000110010000011101101111110111100001110010111100100111100101101011000001110111001011001111000111100000101010110101110101011111110111110101110100000010010001011110100011100010001011111000010001000000111000001000001100111011110000111101011010000111011001110001010011000100001100000000011110000000000011010101000111111001110011111100000100101000111100001101001101111110011001101111110011011111111101111111111000011111100110110001001100100101000011100010100010010111010011100100110110101011000100111011111010010000000011110000100000011110011101101110111111010001101110111001101000001001110000110010101010000100110110101011111110101011101110001000100101111000110010011101111000101000110000110010000000111000001101010010000001111111100010101111001000000111110111100011010101001010110000101111111000101110010001110010111011010110000101100000100010101101110001100011000100010111101100101000101011110001011011010110111000110010010101010010101111000001111110010010010010010000111111101101000010100000101010011101001100101000010110110110111001001010010110101101011110011110011110001110010001010011011111010100000101111001000001101111110010110111000000010101001010110101110111101011001111011101101111101000101100010000111001111011000100011001011100010011111111100010111101010111010001110011100101011000111101001111110010111100100010111000100011101001011100001011101000101011000100110101100101011011110110001000101011111101101110110000010111001011011000100010110100011111010011110101001101010011111101011111010000111110001011100010001101100011111100000011101100001010000010110010111000111111011111110000100101011011100000011010011100110101111011000000111011001010011110010010111100110100110010000010100011110001111100001001010011100101000110110101111010110110100010111000101111100011001100111000110011110110100110001100010110001001101001111001000011000011000010011101101100111100110111000101111100111001010011001100000100001100010000011110011000111000000101110101011111001000101101111100111110100001111100100100000100011010010110000011001100010101110111011101110101101110010011011000101111001001010001110010101010110100100111101111100111101110010101100101011110110010000110010110001110001110011000100001101110111000000000100110010001001111111000010110010111100010000100100001001001100001100010111111100111001001010101100000111000010001001100011100100010011010111101000011010111000101001101011101101010101011101000001010011110010110001001011010001101011100011011011010110101010110001110011000001110111110001111100001111110111001011010110011100101010001111100000011001101110100110101000110011011001011001010110010010110111110010101011011110011001111110100111101100000111010011011001010001001100001010101000000110001011110001010111001000110001010111101110101101101101100111010101010010101110001011100010110111111010001001111000001001110110111100011010111000111110111000100010110010111111111001001001101011000111000011001001110100101011101011111101010100011100100111001011111010000100110110110011000110001100101010111111000100101101001110011001111110010101101110110000110110101011010011110000001010001110000010110100000100011110011100000000000110010110101110101001111100100011000110111100000100110000010000000001101111101001011001100011110100110111100010101111110000010011001110101100011011111110010010111011000001111101100101010101011100000111001001011101010000001000110001001101000101100101110110010100001011001001000001001001111111001100101001000111010100100001000110011010110000010010010000110101101100111001000110001010010011010110100110001011010011001110111101011110110000011101000110000010000001110010001011000000101111001110100011011111001100010000010011111101010000000011011101100110110111011011001011110100101010101101110011000010110011100110100000100111110010011101001011111101100110100101011010001011110000011110011010101011110000000100000000111000000011111010000111111010011000101010100111110010100000001000010001001110101010011010110000100001110101101110011010111101011000010011001100000110011011111000001100000111110011100110111000010011111111010110000000001000110110011001110001011011110001101001010011010000000001110111111110001111101001010001000100111111110001011110100111010000000011000011111101111100000100010010010010111010000101111110011000000011111110111111111111000101111010011010110101000111100111001001111111111001001101011000000101010001000001010101111010100100101101101110011110111110010100110101111010101110000000110011000100011111111111100001001011010110011101101101010110011101111111110100110110011000111001110000111010110010100010101000110011000011001001010011010011101010010100000001110111010000111110110011101000110001000010100010001100010100101000011001100011110101111100111000001100100010111111111010101110110100011010010101010010101011000000101000100011000111010011000001110110111111010111000001010000111111111001000110100011110000011000001001010110110100110101100000010110111010010001000111111101010111100010101110101011000000011001010101000100001010011000000110011100100111111111000100001010010100000111001000000111101100111010000111111011111110111100100001101000000111011010100110101111101011011011111110010100110110000000001011011111100011111011011011111110111011110001111101000011010001100111000001101110000110110001111110110010100100011011000110011100110110100000010000101001010110101111101010110100011100101000000110111000000001000101011100011111011100001110111001010110010101011100001011000011100111001001101111000001101100011000000110111011111011001001010000111100010110010111111110100011110011111100011111111011111111001101011011001; 
		
	end
end

endmodule
