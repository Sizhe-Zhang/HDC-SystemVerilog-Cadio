module random_index_block(
	letterReady,
	inputLetter,
	textDone,
	textVector,
	clk,
	rst
);
parameter N = 10000;
parameter PRECISION_RI = 31;
parameter MAXLETTERS = 10;

input [4 : 0] inputLetter;
output reg [N-1 : 0] textVector;
input clk;
input rst;
input textDone;
input letterReady;

int j, seed;
reg [N-1 : 0] letterVector;
reg [N-1 : 0] letter_1;
reg [N-1 : 0] letter_2;
reg [N-1 : 0] letter_3;
reg [N-1 : 0] letter_4;
reg [N-1 : 0] letter_5;
reg [N-1 : 0] letter_6;
reg [N-1 : 0] letter_7;
reg [N-1 : 0] letter_8;
reg [N-1 : 0] letter_9;
reg [N-1 : 0] letter_10;
reg [N-1 : 0] letter_11;
reg [N-1 : 0] letter_12;
reg [N-1 : 0] letter_13;
reg [N-1 : 0] letter_14;
reg [N-1 : 0] letter_15;
reg [N-1 : 0] letter_16;
reg [N-1 : 0] letter_17;
reg [N-1 : 0] letter_18;
reg [N-1 : 0] letter_19;
reg [N-1 : 0] letter_20;
reg [N-1 : 0] letter_21;
reg [N-1 : 0] letter_22;
reg [N-1 : 0] letter_23;
reg [PRECISION_RI-1 : 0] posCounter [N-1 : 0];
reg [31 : 0] counter;
reg [N-1 : 0] letterEncoding [MAXLETTERS-1 : 0];
reg [2 : 0] state;
wire [N-1 : 0] tetagramVector;


// Shift registers and compute tetagram
always @(posedge clk) begin
	if (!rst) begin	
		for (j = 0; j < N; j = j + 1) begin
			posCounter[j] <= 0;
		end
		letter_1 <= 0;
		letter_2 <= 0;
		letter_3 <= 0;
		letter_4 <= 0;
		letter_5 <= 0;
		letter_6 <= 0;
		letter_7 <= 0;
		letter_8 <= 0;
		letter_9 <= 0;
		letter_10 <= 0;
		letter_11 <= 0;
		letter_12 <= 0;
		letter_13 <= 0;
		letter_14 <= 0;
		letter_15 <= 0;
		letter_16 <= 0;
		letter_17 <= 0;
		letter_18 <= 0;
		letter_19 <= 0;	
		letter_20 <= 0;
		letter_21 <= 0;
		letter_22 <= 0;
		letter_23 <= 0;	
		state <= 0;
		counter <= 0;
	end
	else 
		if (letterReady) begin
			
			letter_23 <= letterVector;
				
			letter_22[N-1] <= letter_23[0]; 
			letter_22[N-2 : 0] <= letter_23[N-1 : 1];		
			
			letter_21[N-1] <= letter_22[0]; 
			letter_21[N-2 : 0] <= letter_22[N-1 : 1];


				
			letter_20[N-1] <= letter_21[0]; 
			letter_20[N-2 : 0] <= letter_21[N-1 : 1];		
			
			letter_19[N-1] <= letter_20[0]; 
			letter_19[N-2 : 0] <= letter_20[N-1 : 1];	

			letter_18[N-1] <= letter_19[0]; 
			letter_18[N-2 : 0] <= letter_19[N-1 : 1];	

			letter_17[N-1] <= letter_18[0]; 
			letter_17[N-2 : 0] <= letter_18[N-1 : 1];		
			
			letter_16[N-1] <= letter_17[0]; 
			letter_16[N-2 : 0] <= letter_17[N-1 : 1];	

			letter_15[N-1] <= letter_16[0]; 
			letter_15[N-2 : 0] <= letter_16[N-1 : 1];	

			letter_14[N-1] <= letter_15[0]; 
			letter_14[N-2 : 0] <= letter_15[N-1 : 1];	

			letter_13[N-1] <= letter_14[0]; 
			letter_13[N-2 : 0] <= letter_14[N-1 : 1];		

			letter_12[N-1] <= letter_13[0]; 
			letter_12[N-2 : 0] <= letter_13[N-1 : 1];	

			letter_11[N-1] <= letter_12[0]; 
			letter_11[N-2 : 0] <= letter_12[N-1 : 1];		

			letter_10[N-1] <= letter_11[0]; 
			letter_10[N-2 : 0] <= letter_11[N-1 : 1];	

			letter_9[N-1] <= letter_10[0]; 
			letter_9[N-2 : 0] <= letter_10[N-1 : 1];		

			letter_8[N-1] <= letter_9[0]; 
			letter_8[N-2 : 0] <= letter_9[N-1 : 1];		

			letter_7[N-1] <= letter_8[0]; 
			letter_7[N-2 : 0] <= letter_8[N-1 : 1];	

			letter_6[N-1] <= letter_7[0]; 
			letter_6[N-2 : 0] <= letter_7[N-1 : 1];	

			letter_5[N-1] <= letter_6[0]; 
			letter_5[N-2 : 0] <= letter_6[N-1 : 1];	

			letter_4[N-1] <= letter_5[0]; 
			letter_4[N-2 : 0] <= letter_5[N-1 : 1];	

			letter_3[N-1] <= letter_4[0]; 
			letter_3[N-2 : 0] <= letter_4[N-1 : 1];	

			letter_2[N-1] <= letter_3[0]; 
			letter_2[N-2 : 0] <= letter_3[N-1 : 1];	

			letter_1[N-1] <= letter_2[0]; 
			letter_1[N-2 : 0] <= letter_2[N-1 : 1];	

		
			if (state < 23)
				state <= state + 1;
			else begin
				counter <= counter + 1;			
				for (j = 0; j < N; j = j + 1) 
					if (tetagramVector [j] == 1'b1)
						posCounter[j] <= posCounter[j] + 1;	
			
			end
		end
end

assign tetagramVector = letter_23 ^ letter_22 ^ letter_21^ letter_20 ^ letter_19^ letter_18 ^ letter_17^ letter_16 ^ letter_15^ letter_14 ^ letter_13^ letter_12 ^ letter_11^ letter_10 ^ letter_9^letter_8 ^ letter_7^ letter_6 ^ letter_5^ letter_4 ^ letter_3^ letter_2 ^ letter_1;

// Do thresholding based on counter values
always @(posedge clk) begin
	if (!rst)
		textVector <= 0;
	else
		if (textDone) begin 		
			for (j = 0; j < N; j = j + 1) begin
				if (posCounter[j] > (counter >> 1))
					textVector[j] <= 1;
				else
					textVector[j] <= 0;
			end
		end
end

//initial begin
always @(posedge clk) begin
	if (!rst) begin	
		letterEncoding[ 0] <=10000'd0;
		letterEncoding[ 1] <=10000'd0;
		letterEncoding[ 2] <=10000'd0;
		letterEncoding[ 3] <=10000'd0;
		letterEncoding[ 4] <=10000'd0;
		letterEncoding[ 5] <=10000'd0;
		letterEncoding[ 6] <=10000'd0;
		letterEncoding[ 7] <=10000'd0;
		letterEncoding[ 8] <=10000'd0;
		letterEncoding[ 9] <=10000'd0;

	end
	else begin
		letterEncoding[ 0] <=10000'b1100101100111001011111010110101010110110110101011111101001001110010001101011000001111100001100011010001101110001001111001110000110001110110010111010011001110000010111110001111000011001000001001111001010010010000100000011101010111010111100100011001001001111111101000100110100110110101000101101101110100000100111100011010110000000101001011110010111000110011000111111010001001100100010111010101101111011100000001001011011110100000001100111010011001011110011101110010100111001110001101000000000010111110101010011000000000100011110011001000100010100101100110100110110111011011110011000011100100001111011001011100100101011100001011010111100001010110000101000011001101010111100101010111011101100101001111100111110101110110001011101011010101100011001101011000110111001011110010000111010101011111010000110101010110000101011010000101000000100111101111011001000000000100011100011100101001100110101011100100010101101100011101100101010011011000101101000111011100010000010001000110000100101110010000101011110110101111010011000001111011100010000011111000110100111110111001110001110011111011111010000001001101011110111011101000111110110110011011111110011011110110110001001010101001100110110100010011101011111110010110001010000101100110010101011011101101101010111011111001111110011110110101010100101011110001011100100110000111111001011110100011111100010011011110101111110110101001010110011101001001110111100111001110111000101110000111001110110000010000111111011100111000111011010111110000111111110010110111111010111001110000000100000111010111111110100100101000101110011010100100000111111010010000101101110111110001110100010100001011110000011010011100111010100111111111010010110000011101110000100001011110010101010011100111110110000110100110110001010111111100011100101111110010110001101000100000010101001101110000010100001101010000100111100111110010010100011010101000100010110000001111100010101111010000011111100100101000010111011111111000001111101010111001111101010011111111100011001100111010110001011000111111110001011100011000010010010100101110010111001111011111100100000011110101111111010001101001000001001101000001011110110010101110010010001001001001111100101110011001000100010000010111110100001111101100101011011110000011100111011111001101001101000001100011011110101010010111110110110110101100010100111111011110111101011110001010101001101010000000101011111100111100011001010111010100111101100010000110101111101010000101011111011001101111000011001100011111001001000011110010110001010101100111100010000100011000101111001100100110001000011011101111110110001011111001010111100110101000010101000100011100001100000000100000001000111001000011001000111010101100111011011101010110011101010010001000100101110010100110001001001001100001101111111110000011111010001110101010101010111100100101110111011111010010110110010011001111100010000011000010011010000011110110000010001110101111011000101111010010011101100101101010011010001011111000010001001010111001110100011010111111111001010100001100100000000000101011110001001001000001011001101110101000010010111101011110010000110011100100001011010010001100001010011000000000110000110011101110011011110111100100100101111010000000100101000011101111111101100001001000000111010011100001001110000011000000010110001000110010111101111111001000100100100010111100101000000101111000001111001000000100101111000100000000101111010010110110010000011100001000101000110111111010110101101010011001100110100001000100101001011010011001111010100001101111100001010011110000011000111110100000101011100100110011001111001111010100011110011100000010011001010111111011000001001011110010011010000111011010011001000100101000100010001101101111010001111010110111011111000001100101110000111100010010000101011011100011001000000001010100001000001011001110111001110111010101000100001110110110110111101010010000000000111001100001011011001111101011100101010110100011010100000101000100100100111101000110101100000001011001000001111100101100111110100100101010010010111000100101100001100101110010111100011010001010000111011111010001111011011010000101111000001100000100000101001101000110000010100001100000111111010001111011101000110100101111111000110101001000111010000001000110110101001100001101110101010110101101111000101100110101111001110101010100011101101000011010110101010101111110011010101110110101010000100001010110101011100100011110111011110001110011001110111110110111001111001000110010000110100010011010001011000100010000001100111111110111010001111010010000111001111110001000110010001100100111110001111010011110000010010110010101011110000011001001110110011100000010101000011000111000000000010100010100100010110010010100011110110000010000100110111101110111011111101110001100001111010110100101101101111000101001110101111000111110111010110110001101000110111101001000011011111011111010011101001010111110001101111011100101001010101010001001100110111011000001011111100110000101000011101110101011001010010000101111100101110010100000110001111110111111100001010101000100111111010101101000101000011101110011100100011110001110001110111100110100100001101101011100101000011000000001111011101010100101000110000110100000111000001111100010011111110010001010010001111101010010000011010111110100110011001110110011011111011100001111111111010010000100001000000110010011101101100001010010101010010101010101100010111111101000101111101111101010011101010011000100101110101111110100100111001101111100110100010000000011101001010001010110110000010010100110000110101110010010000101010011100100100110011101110111011000000100000000011111001011011001001110111000111101111100101011010011100010100110011110101000101011101011011000111100111110001001001011111111110010100010110111111011000101010001010001000100101100011101111101000001110000101110111000001110110100001110101000000100101100100010001101100001011001110000110011100101110000101110111101100110111101111111010110111010111011101110011001010010111101111101001110101000110011110000011010000001000110011110010011101100111001011000110010001011111111111010011111110110000000000111111010000010000101011011111010101110101110001111101111001101010011100100100001000001111100001000011101100001100000000011111000001111010010011010001110011110100101001100011010010000000000011000111011010100000110000001000101011011101101110111011110001101010000000001011000110100001111111000111110001011010011111111000000111101111001110001101100110010101010001011111011001110010110100001111101100011011000010010001100000111010010101111011100010001110011000100101110110111000011111110101010010011011001001001110000100000100101011011100000110010001000110101011000000100101010111011011110100110100101111100000111011001011010001110110000111010011101011010100011000001001011000100001001101010001101110101011101010000010001010100110111100100011111110000111011011101101101101101111101110110111000011001111011110100100110110100100001001111011100001100101101000101000111110011010110000010100010010001010010110001011010001101010010101110000011110110100001001010000110010001110001000011110000000110000010111001011100000011101011101000000101100101110110101110011011001100011001001011100110000101011111111001111111010001111110100001001101101110111001111111011010101000011110111001001000101011100000000111101100111011011110100100111000101000101110101110010010111001101011110000011000010001100011101001011100101111001001010010000100110010000001000110100101011100101001000000110111111001001011000000011110001001010111111111100101111001100011100010111000001010001101111011001110110000001000001000000010011101011001010001011010111100011000111001101110000101011000010101101100000011001110101010010011001101010000011000000100011010001010000010001001100100000100001100100010101110101000100110100001000101100111101000000100100011111010110001010100111001101010111001000000101101110100000010010011101010100000101001101001011100001010001000100111110100010010000101010010011111011100110101111101110001000010000010101000111101111010110100001000111000010100011011111001111011110111011010110101100000110100011000000111010001000111110110001001101011001010110101110000100010110011101010111100100001011000010101011111111011001111111010000000001000111001100101011000000000010100100010000110011101110000110101010111111100101000011011100100111000101110001001100000011001101000110110100101010000001011001111001100111001100001101010100111001110110100001001001001110011101001001101101001111101111000010110101111000000110011111000011111000100010000101010000100011100111010010011110110100001110011101010010010100111110011000111000101110010000110110000110111000110110100100111001110010110010000000000010001111000100110111101011100011011101000001001010100010101001100101100001001100100110111111111110000001110101101011011001101001110110100101000000111011101110011010000010100010111000110101001011100111111111010011111011010000100011100010001011111111000001001101110100010101010001011110110011011010011001100100100111111100010100000001111110111111001101011010010000110000111011100001001001011001111011011011100011001010111001111001110001100101010111100001010000000001110100010011000111100110100110110001110110011000100110001011111111011100101010110100010101010110001100111110111111111000100101110001100110100100011010000000101000101110001000101011011010000001011001100010101111101011110010000110001101101100000101110101111001100011111011000010111010000001100001101100001000100000011100011000101111001110100101110001100111110101010000100111111111111010110101010101011111011111110111111101010110110010000101001000000000000001101111010111111101000010111010110001001000010101010010011101100110101011001111010011010110011110100101110000111100001011000110100110110111001101001010000000001110010000101010011101001111100110101101001011110001101011101101010110100010011110111111000110100011111001011111100110001011110010011010001110001111001000100110010010111011111001011100101101110000001101111111010111001011010010010011011001110000100100110000001111010001010000000000110110110101010011011100010001000100000011110010010010010101010101110010011001100110111111000000010111; 
		letterEncoding[ 1] <=10000'b1100101100111001011111010110111010110110110101111111101001001110010001101011000001111100001100011010001101111001001111001110000110001110110010111010011001110000010111110011111000011001000001001111001010010010001101000011001010111011111100100011001001000111011101000000110100110110101000101101101110100000100111100011011110000100101001010110010111000110011000111110010001001100100010101010101101111011100000001001011011100100000001100111010011011011110011101110010100111001110001111100000000010111100101010011000000000100011110111001001100010100101100110100110110111011011110011000011100100001111011001011100100101011100001011010111100001011110000101000011001101010111100101010111011101100101001111100111110100110110001011101011010101100001001101011000110111001011000011000111010101011111010000110101010110000101011010000101001000100111101111011001000000000100010100011100111001100110100011100100010101101100011101100101010011011000101101000111011100010000110001000110100100101110010000101111111110101111010011000001111011100010000011111100110100111110111001111000110011111011011010000001001101011110111011101010111100110110011011111110011110110110110001001010111101100110110100010011101011011110010010001010100101100110011101011011101101100011111011111001110110011110110101010100101110110001011000100100000111111001011110100011111100010011111110101111110110101001011110011101001011110101100011001110111000101110000111001000110000010000111111011100111000111011010111110000111111111010111111111010111001110000000100000111010011111110100100101000001110011010100100011111111010010000101101110111110001110000010100001011110100011010001100101010100110111111010010110000011101100000100001011110010101010011000111110111000110100110111001010111101100011100101111110011110001111000100000010101001101110000010100001101010000100111100111110010010100001011101000100010110000000111100010101101010000011111100100101000010110011111110000010101101000111001111101010001111111001011001100111010110001011100111111110001011100011000010010010100101110000111001110011111100100000011110101111111010001101001000001001101000001011110110010101110010010001001011001111101101110011001000100010000010110110100001111101100101010011110101011100111011111001101001101000001100011011110101010010111110110110010101100010100111111011110101101011110001010001011101010000000101011111100111100011001010111010100111101100010000010101111101010000101011111001001101111000011001100011111001001000111110000110001010101100111100010000100011000101111001100100110001000011011101111110110001011111001010111100010101001010101000100011100001100000000100000001000111001000011011000111010111100111111011001000110011101010010001100100101110010100110001001001001100001101011111111100011111010001011001010101010111100100101010111011111010110110110010011001111110010000011010010001000000011110110000010001110101111011000101101010010011101100101101010011010001111111000010001001010111001110100011010111111111101010100001100100000000000101011110001001001000001011001101110101000010010111101011110010000110011100100001010010010101110001010011000000000110000100011101110011011110111100100100001111010000001100101000011101111111101100000100000100111110011111001001110001011001000110010000000110010111101111111001000100010100010111100111000000101111000001111100100000100101111010100000010101111010010110110010000011100001000101000100111111010101101101010011000100111100001000100101001011010011000111010100001101010100001010011110000011100111110100000101011100110110011001111001111010100011110011100000010111001010111101011000001001011110010011010000111011010011001000100101000100010001101101111010001011000111011011111010001100101110000111100010010000101011011100011000000000001010000001000001011001110111001110111110101000100001110110110110111101011010001000000111001100001011011001111101011100101010110100011010100000101010100101100111101000110101000000011011001000000110100101100111110100000101010010010111000000101100001101101110011111100010110101010000111011111010001111011011010000101111000001100000100000101001101000110000000100001100000111110000001111011101000110100101111111000110101001000111010001001000110110101101110001101110101010110000111111000100100110101110011110101010100011101101010011010110101010101111110011010101110110101010001100001010110101011100100011110111011100001110011001110111100110111001111001000110010000110100010011010001111000100010100011100111101110011000001101011010000111001111110001000110010001100100011110001111010010110000010010010010101011110000011001001110110001100000010101000011000111000001000011100010100100010110010010110011110110000010000000100111101110111011111101100001100001111010110100101101111111000101001110101111000111110111010110110001101010110111101101000001010111011011010011101101110111110101101111011000101001010101010000000100110111011000001011110001110000101000011101100101011001010110000101111100101110010101000110001111110111111100001010101000100111111011101101000101000011101110011000100111010001110001110101100110100100001101101011101101000011000000001111011101010100101000110000100100000111000000111100010011111110010001010010001111101010010000011010111110100110011101110110011011111011100001111101111000010000100001000100100000001100101100001010010101010010101010100100010111111101000101111101111101010011101010011000110101110101111110100100111011101111100111100010000000011101001010001110110110000010001100110100110101110010010000101010011100100100110011101110111000000000100000000111111001011011001001010110000111101111100100011010111100010100111011110101000100011101011011000111001111110001001001001111111110010100010110111111011000101011001110001000100101100011101111101000001110000101110111000001110110100001110101001000100101000100010001101100101010001110000110011100101110000101110111101100110111000111111010110011010111011101110011001011010111101111101001110101000110011110000011010000001000110011100010001101100111001011000110010000011111111111010011111110110000000000111111010000110000101011011111010101110101110001111100111001101011011100100100001000001111100011100011101100000100000000011011000001111010010011010001110010110100101001100111010010000000000011100111011010100000010000001000101011011101101110111011110001101010000000001011000110100101111111000111110001011010011111111000000111101111001110001101100110010101010001011111011001110011110100001111101101011011000010010001100000111110010101111011100010001110001000100101110110111000011111110101010010011011001001011110000100000100101011011100000110010001001110101011000000100101000011011011110100100100101111100000011011001011010001011110100111010011101011010100011000001001001000100001001101010001101110101011101010000010001010100110111100100011111110000111011011101101101101101111101110111110100111001110011110100100110110100000101001111011100001100101101000101000111110111010110000010100010010001010010110001011010001101010010101110010011110110100001001010000110010001110001000011110000000110000010111001011100100011101011101000000101100101110110101110011011001100011001001011100110000101011111111001111110010001111110100001010101101110110001111111001010101000011110011001001000101011100000001111101100111011001110101100111000101000101110101010010010111001101011110000011001010001100011101001011100101111011001010010000100110010000001000110100101011100101001000000110111111001001010100000011110001001010111111111100101111001100111100010111000001010001101111001001110111000001010101000000010011101011001010001010010111110011000111001101110000101011000010101101100000011001110101010010011001101010000011000000100011110011010000010001001100100000100001100100010101111101100100110110011011101100111101000000100100011111010110001010100011001101011111001000000101101110100001010010111001010100000101001101001001100001010001000100111110100010010000101010010011111011110110101111101110001000010101010101010111101111010110100001000111000010100011011111001101011110111011010000101100000110100011010000111010001000111110110001001111011001010110001110000001010110011101000111100101001011010000101011111001011001111111000000000001001111001100101011000000000010100100011000110011101110000110101010011111100101000001001100100111000001110001001100000011001111000110110100101010000001111001011001101011001100001101010100111001110110100011001001001110011101000001101101001011101111000010110101111000000110011111000011111000100010010101010000101011100111011010011110110110001110011101010010010100010111011010111000111110010100110110000110111000110110100100111001110000110110000000000010001111001100110111101011100001111101000001001010100010111001100101100000000100100110111111111110000001110101101010011001101001110110100101000000111011101110011000100010100010111000110101001011100111111111010011101011010000110011100010001011111111000001001101110100010101010001011110110011011010011000100100100110111100010100000001111110111011001101111110010000110000111011100001001001011001011011010011100011001010111101111001110001100101010110000001010010000001110100010011000111100110100110110001110110011000100110001011111111011100111010110100010101010110001100111110111111111000100101110001100110100100011010100010101000100110001000101011101010000001011001100011101111101010110010000100101101101100010001110101111001100011111011000010011010000001100001101100001010100000011100011000101111001111100101110001100111110111010000101101101101111010110001010101011111001111110111111101010110110010000101001000001000000001101111110111111101100111111010111001001000010101010010010101100010101011011111010011010110011110100101010000111110001011000110100110100111101101001110000000001100010000101011011101001111100110101101011011110001101011101101011100100010011110111111000110000011111001011111100110001011110010011010001110001111001000110110011010111010111101011100101101100000001101111111010111001010010010011011111001100100100100010000001111000001010000010000111110110101010011011100010001110110000011111010010010010101010101100010011001100101111111001000010111; 
		letterEncoding[ 2] <=10000'b1100101100111001011111010110111010110110110101111110101001001111010001101010000001111100001100011010001101111001001111101010000110001110110010111010010001110000010111110011111000011101000001101111001010010010001101000011000011111011111100100111001001000111011101010000100100110110101000101101101110100000100111110011011110000100101000110010000111000110011000011110010001001100100010111010101101111011100100001001011011100100000001100111010011011011110111101110010000101001110001111100001000010111100101010011000000000100011110111001001100010100101100110100110110111011011110011000010100100001111011000011100100110011100001010010111100001011010000101000010001101010011100100010111011101100101001111100111010000110110001011101011010101100011001101011010110011001011000011000111010101011011011000110101010110000101011010000101001000100111101111011001000000000100111100011100001001100110100010100101010001100101011101100101010011010000101101000111001100010100110001000010100100101110010000101111101110101011010011000001011011100010000011111100110110111110111101110000110011111011011010000001011101010110111011101010110100110110011011111110011110110100111001101010111111100110110100010011101011011110010010001010100101100110011101011011101111100011111001111001110111011110110101010000101110110001010000100100000111111001011111101011111110010111111110101111100110101011011110011111101011110101100011001110111000101110000011001000110000010000111111011100011000111011010111110000111111111010110110111010111001100000000100000111010011011010100100101000001110011010100100011111110010010000101101110111110001110000000100001011110100011010101100101010101110111111010010110000011101100000100001011100010101000011000111110111000110100110111001010111001100011100101110110011110001101000100000010101001101110000010100001101010000100111100111110010010100001010101100000010110000000111100010101101010010011111100100101000010110011111110000010101101000111001111101010001111111001011001100111010110001011000111111110001111100011000010000010100111110000011001110111111100100000011010101111111010001101001000001001101000001011110110011101110110010001001011001111101101110011011000100010000110110110000001111101100101010011110001011100111011111001101011101000001100011011010101010010101110100010000101100010100111111011110101101011110001000001011101010000000101011111100111100011011010011010100111100100010100110000111101000000101011111001001101111000011001100011111001001100011110000110001010101101111101010000100011010101111111100100110001000011011101111110110001011111001010111100010100001011101000100011100001100000000100100001000111001000011011000111010111100111111011001000110011101010010001100100101110010100110001001000001100001101011011111000010111010001011001010101011111100110101010111011111011110110110010011001111110110100011010010011000000011110110000010001110101111011000101101010010010101100101101010011010001111111000010001001010111001110100011010111101111101010100001100100000000000101011110001001001000101011001101110111010010010111101011110010000110010100100001010000010101110001010011000000000110000100011101100011011110111101100100001111010001001100101000011101101111101101000100010100111110011111001001110001011001000110000000000110010111101111111001000100001100010110100111000000101111000001111100100000100101111010100000010001111010010110110010000110101001000101000100111111010101101101010011000101111100001000100101001011010111110111010100001101010100001010011110000011100111110100000101011100110110011011111001111000100011100011100000010111001010111101011000001001011110010011010100011011010011001000101001000100010001101101111010101001000111011010111010001100101110000111100010010000101111011100011000000000001010010001000001011001111111001110111110101000100001110110110110111101011010001000000011001100011011010001111101011101101010110100010010100000101010100101100111101000110101000000110010001000000110100101110111110100000001010010010111010000101100001101101100011111100010110101011000111011110110001111011011010000101110010011100000100000101001101000110000000100001100001111111000001111011101000110101101111111000010101001000111010001001000110111001101110001101110101010110000110111000100100110101110011110101000100011101101010011010110101010101111110011000101110110101010001100001011110101001100100011110111011100001110011001110011100110111001111001000111011000110100010010010101111000100010100011100111101110001000001101011010000111001111110001000110010101100100011110001111010010111000000010011010101011110000011001001110110011100000010101000011000011010000000011100110100100010110010010111011110110000011000000100111101110111010011101100001100001111010110100101101111110000101101110101111000111110111010110110001101010110011101101000001010111011011000011101101110011110101101111011000101001010101010000000000110110011000001011110001110000101000011101100101011001110110000101111100101110010101010110001111110111111100001110101010100111111011101111000101000010101010011000100111010001110001110101110110100101001101101011101101000011000100001111011101010100101000110000100100000101000000111100010011111010010001010010001111101010010010011010111110100110011101010110010011111001100001111101111000010000100001000100101000101100101100001010010101010010100010000100010111011101000101111101101101110011101010011000110101110101111110100000111011000111100111100010100000011101001010001110110110010010001100110100010101100010010000101010011100100100110011101110111000000000100000000111111001011011001001010110010111101111100100010010011100010100111011110101000111111101011011000111001111100001001001001111111110010100010110111111011000101110001110001000100101000011101111101000001110000001110111000001110110100001110101001000000001000100010001101100101011001110000100011000101110000101110101101100110111100111111010110011110011011100111011001011010111101011101001110101000110001110000011010000100001110011100010001111100111001011000110010000001011111111010011111110110000000001111111011000110000101011011111010101110101110001111100110001101011010100100100011000101011100011100011101100000101000000011011000001111010011111010001110010110100101101100111010010000000000011100111011110100000010000001000111011011101101110111011110001101010000000011011010110100101111111000111100001011010010111111000000111101111001110001101000110010001011001010111011001110011110100000111100101011011000010010001100000111110000101111011100011001111001000100101110110111000010001110101010010011011001001011110000100001100101011101100001100110001000110101011000000100100000011010011110100100100101111100000011011001111010001011110100111010011101001010100011000000001011000100001001101010001101110101011111010000010001010100110111100100011111110000111011011111101101101101111101110111110100111001110011110100100110110100000100011111011000001100101101000101000111111111010110000010100010010001010010110001011010001101010010101110010011110110100001001010000110010001110001000011110000100110000011111001111000100011101011100000001101100100110110101110011011001100011001101111100110000101011111011000111110011001111111110001000101101110111001111111001010101000011110011001001000101011100000101111101100111011001110101110111000101000101110101010010010110001101011110000111001011001100011101001011101101111011001010010000101110010000011000111100101011100101001000000110011111001101010100000011110001001010111111111110101111001100111000010111000001010001101111001000110111000001010101000000010011101010001010001010010111110011000111001101110000111011010010101101100110011001110101010010111001101010100011000000100011110011010000010000001100100000100001100100010101011101110101110110011011101110111101000000100100011111010110001110100011001101011111001101000101101111100001010110111001010000000101001101001001100001010001000100101111100010010000111110010011011011110110101111101110001000010101010101010101101110110010100001000111000010100011011111001101011110111011010000101100000110000011010000111010001000111110110001001111011001010110001100000001011110011101001111100101001011010000101011111001001001111111000001000001001111001100100011000000000010100100011000110011101110000110101010011110100110000001001100100111000001110011001100000011001111000110110100101010101001111001011001101011001100001101010100011001110110000011001001001110001101000001101101001011101111000010110101111000000110011111000011111000100010010101010000001011100111011010011110110110001110011101010011010100010111011010111000111010010100110110000110111000110100100100111001110000110110000000001010001111001100110111101011100001111101000001001010100010111001110101100000000100100110011111111110000001110101111010011001100001110110100100000000111011110110011000100010101010111000110101001011100111111011010011101011010000110011100010001011111110100000001101110100010101010001011110110011011010011001100101100110110100010100000001111110111011101100111110010000111000111011100001001001010001011010010011100011001010111101110001110001100101010111000001000010100011100100010001000111000110100110110001110110011000100110101011111111011100111000110100010101010110001100111110111111111000100101110001100110100100011010100010101000100110001000101111101011000001001001100011101110101010110010000100101101101100010001110101111001100011111010000110011010000111100001101100001000100000011100011100001111001111100101110001100011110111010000101001101101111010110001010101011111001111111111111101010111111010100101001000011000000001101111111111111101100111111010111001001000010101011010010101100010101011011111010011010110011111100101010000111110001111000010100110100111101101001110000010000100010010101011011101000111100110101101011011110001100010101101011100110000011110111111000110000011111001011111100110001011110010011010001110011111001000110110011010111010111101011000111101100101001101111111011111001110010010011011111001100100100100010000011111000001010000010100111010110101010011011100010001110110000011111010000010010101010101100010011001100101111101001000010111; 
		letterEncoding[ 3] <=10000'b1100101100111000010111010110111010110110110101111110101001001111010011101010001001111100001100011010001101111001001111101010000110001111110010111010010001110000011111111001111001011111000001101111001010010010001100000011000010101011101100100011001001000111011101010000100100111110101000101101101110100000100111100011011110000100101000110110000111100110011000011110010001001101100000111010101101111011100110001001011011100100000001100111010011011011110101101100010000101011110001111100001100010111100111010011000000000100011110111001000100010100101100110100110110111011111110011100010100100001111001000011100100110011100001010100101100001011010000101000010001101010011100100010111011001100101001111100111010000110110000011100011010101100011001101001010110011011011000011000111010101011011011000110101000110000111011010000101001000100111101111011001000000000100111100011100001011100110100000100101010011100100011101110101010011010000101101000111001100010110110001000010110100101110010000101111101100101001010111000011011011100010000011111100110110111010110101110000110011111011011010000001011101010110111011101010110100110110011011111110111110110100011001101010101111100100110100010011101011011110010010001010100101100110011101011011101111100010111001111001110111011110110101010000101110110000010000100110000111111001011111101011111010010111101110101011101110101010011101011111101011110101101011001100111000101110000011001000110000110000011111011100011000111011010111110000111111111010110110111010111001100000000100000111000011011010100100101000001110011010100100011111110010010000101101110101110101110000000100001011110100011000101100101010101110111111010010110000001101100000100001011100010101000010000111110111000110100110111001010111001101011110101110110001110001001000100000010101001101111010010000001101010100100111101111110010010100101110101100000010110000000111100010101101110010011011100100101000010110011111110000010101101000111001111101010001011111001011001100111010110001011000111111110001111100011000010000010100111110000011001110111111100100000011010101111111010001001101000001001111000000011110110011101110110010001001011000111101101110011111000100010000010110110000101111101000101000011110001011101001011111001101001100100001110011011010001010010101111110010000101100010100010111011110101101001110001000001011101010000000101011111000111100011001010011010100101100100010000110000111101000000001011111001001101111001011001101011111001001100011110000110001010101101111101010100100011010101111111100101110001001011011111111110110001011111001011111100010100001011101000100011100001100100000100100001000111001000011011000111010111100111011011001010110011101010010001100110101110110100110001001010001100011101011011110000010111110001011001010101011111100110111010111011111011110110110010011001111110100100011010010011000000101110110001010001110100111011000101101010010010111100101101010011010001111111000010001001000111101110100011010111101111101010100001100100000000000101011110101001001000101011001101110111010010010111101011110010000110010100100001010000010101110011010011000000000110001100011101100011001110111101100100001011011001001000101000011101101111101101000101010100111100010111001011010001011001000110000000000110010111101111111001000100001101010110100111000000101111000000111100100100100101101010100000010000111010010110110010000110101001000101000100111111010101101101010011000100111110001000100101111010010111110111010100001101010100001110011100010011000111110100000101011100110110011011111001111000100011100011100001011101001010111101011000001101011110010011010100011011010011001000101001000100010001101101111010101001000101011010111010001100101110000111100110010000100011011100011000000000001010010001000001011001111111001110111111101000100001110110110110111111011000000000000001001110011011010001111101001101101000110100010010100100101010100101100111101000010101000000110010001000000110100101100111110100000001010010010011010000101100001101101100011110100010110101011000111011100111001111011011010000101110011011100000100000101001111000110000100100001100001111111000001111011101010110101101011111000010101001100111010011001000111111001101110001101110111010110000110111000100100111101100011010101000110011101101000011010110001010101111110011000101110110101010001100001001110101001100100010110111011100001110011101110001110110111001111001000111011000110100010010010101111000100010100011100111101110001000001101011010000111001111110001001110010101100100011110001111010110110000000010010010101011110000011001001110110011100000010101100011000011010100000011010110100100010110010010111011110110000011000000100111101111111010011101100001100001111010110100101100111110000101111110111111000111110111010110110001101010110111101101000001010101111010000011001101111011110000101111011000101001010101010010100000110111011000001011110001110000101000011101100101011001110110000101111100101110010101011110001111110111111100011110100010100111111011101111000101001010101010011000100111011001110001110101110001100101001101101011101101000011000100001111011101010100101010110000100100000101000000111110000011101010110001010010001111101010010110011010111110100110011100010110010011111001100001111101110000010010100001000100101010101100101100001010010101010010100110000100010111011101100111111101101101110011101010010000111101110100111110100000111010000111101110100010100010011101011010001110110110010011000110110100010101100010010010101010011101100100110011101100111000100000100000100111111001011011000001010110010111001011100100010010011100010100111011110101000111111101001011000111101111100001001001001111110110010100010111111110011000101100001111001000100101000011101111101001001110000001110111000001110110100001110101001000100001000100000001101100101001011110000100011000101110000101010101101100110111100111111010110010110011011100111111001011010111101011101001110101000110001010000011010000100001110001000010101110100111001011000110010000001010010111010011111010110000000001111111011000110000101011011101110101110101110001110100110001101011010000100100011000101011100011100010101100000101000000011011000001111010011110010001111000110100101001100010010010000000000011100111011110100000010000001000111011011101101110111011110101101010000000011011011110100101111111000111100001011010010111111001000111001111001110001001000100010001001001000111011001110111110100000111100101011011000010010001100010110110000101111011110011101111001000100111111110111000010001110101010010011011001011011110010100001100101011101100001110110101000110101011000000100101000011010011110100100100101111100000001011001111010001011110100111010011101001011100011001100001011010100001001101010001101110101011111010000110001010100110011100100011011110000111011111111101101101101111101110111110100111001110011110110101110110100000100011111011000001000101101000101000111111111010110000010100010010001010000110001011010001101010010101110010011110110100001001010000110110001110001000011110000100110001011101001011000100011101011101000001101100100010110101110011011001100011001101101100110000101011111011000111110011001111111110001000101101110111000111111001010101000011110011001001000101011100000101111101100111011001110100110111000101100101110101010010010110001101011110000111001011001100011101001011101101110000001010011000101110010000011000111100101011100101001001000110011111001101010110000011110001001010111011111110101111001100111000010111010000010001101111001000110111000011010111000000010011101010001010000010010111110011000110001101110000011011010110101101100110011001110100010010111001101010100011000001100011110001010000010010001100100000100001100101010111011101110101110110011001101110111101000000000110011011010110001110100011101111011111001101000101101111100001011110111001010000000101011101001001100001010011000100101110101010010001111110010011011011110110101111101100001000010101010101010101100010110010100001100111000011100011011111001101110110111011010000101100101110000011010000111010011000111100110001001111011001010110001100000011111111011101001111101101001011010000101011111001001001011111000001000001001111101100100011000000000010100100011000110011101110001110101010011110100110000001001100100011001001110011011100000011001111000110110100101010001001111001011001101010001100001101010100011001110110000011011001101110011101000001100001001011101111000010110111111000100110011111000011111100100010010101010000001011100111011010011110110110001110011101010011010100010110011010111000111010010100110110000110111000110000100100110001110000111110011000001010001111001100110111001011100001110101001001001010100010101001110101100000000110100110011111111110000001110101111010011001101001110100100100000000111011000110011010100010101010111000110101001011100011111011010011101010010000110011100011001011111110100000001101110100010101010101011110110011011010011001100101100110110100010100000001110110011011101100111110010000111000111011100001001001010001011010010011100011001010111101110000110001100101010111000001000010000011100100010001000111000010100110010001110110011000100110101011111011011101111000110100010101011110001101111110110110011000100001110001100110100100011010100010000000100110001000101111101010000011001001100011101110101010110010000100101101101100010001110101111001100001111010000010011010000111100001101100001000101000011100011100001111101111111001110001100011110111110000101001101101111010110101001111011111001111111111111101010111111010110101001000011000000001101111111111111101100111101010111001001000010101011000010101100010101011011111010011011110011111100101010010111110000111000010100110100111101101001110000010000001010010101011011101000101100111101100011010110001100010101101011100110000011110111111000110000011111001011111100111001011110010011010001100111111001000110110011010111010111101011000111101100101000101111111011111001110110010010011111001100010100000000001011111000001000000010100111000110101010011011100010001110110001111111010000010010101010101100010111101100101111100011000010111; 
		letterEncoding[ 4] <=10000'b1100101100111000010111010110111010110110110001111110101001001111110011101011001001111100001000011010001101011001001111101010100110001111111010110010010000110000111111111001111001011111000001101111001010010010001100000011000010101011101101110011001001000111011101010000100100111110001000101001101110100000100101100011011010000100101000110110000111100110011000011110010001001101100001111010101101111011100110001000011011100100000001100111010001111011100101101100010000111011100001111100001100010101100011010011000110000100111110111001000100010100101100010100100110111011111110010101010100101001111001000011101100110001100011010101101100011011010000101000010001101010111100100000111011011000101001111100111010000110110000001000011010101100011001101001110110011111011000011000111010101011011111000100101000110010111011010000101001000100111101111011001000100000100111100011100001011100110100000100101010011100100001101110101010011010000101101000011001100010110110001000010110100101110010000101111101100101001010111100011011011100010000011111100110110111010110101110000110011101011011010100001011101000110111011101010110000110110011011111110111110110100011101101010101111100100110100110011101011011110000010100010100101100110011101011001101111100010101000111001110111011110110101010000101110110000010000100110000101111001011111101011111010010110101110101111101110101010011101011111101010111101101011001100111000101110000011001000110000111000011111011100011000111011010110110000111111111010110100111011111001100000000100000111000011001011100000101000001110011011100100011111110010010000101101110101010101110000000100001011111100011000101100101010001110111111010010110000000101100000100001011100010101001110000111110111000110100111111001010111001101001111101110110001110001001100100000010101001101111010011000001101010110100111101111110110010110101100101101000010110000000111100010101101110010001011101100101000011110011011110001010101101100111001111101011001011011001111001100111010110001011000111111110000110100011000010000010101111110000011100110111111000100000011000101111111000001001101000001001111000000011100110011101110110010001001011000111101101111011110010110010000010010110000101111101000001000011110001011101001011111001101001110100001110011011010001010010101100110010000101100110100000111001110001101001110001000001011101010000000101011011000111100011001010011010100101100100010000010000111101000000001011111001001111111001011001101011111000001101011100000110101010001101111101010100100011000101111111100101111001001011011001111110110001011011101011111000010100001011101000100011100011100100100110100001100111001000011011000111010111110111011011001010110011101010010000100110001110110100110001001010001100010001011011110000000111110001011001011101011111100110111010111011111011110110110010011101011110100100011000010011001000101110110001010001010000111011000101101010010010111100101101010011010001111111000010001001000101101110110011010111101111101010100101100000000100100101011110101001001100101011000101010111010010010111101001010010000110010100100001110000010101110011010011000000000110001100010101100011001110111001100101001011011101001000101000010101101111101111000101010100111100001111100011010001011000000110000000000110010111001111111001000100001101010110100111000000101111000000111100100100011101101000100000010000111010010110110010000110101001000101100100111111010101101101010011000100101110001000100101101010010101011111010100001101010100001110011100010011000111100100000101011100110010011011111001111000100011100011101001010101000010111101011000000101011110010011010100011011011010000000101001000100010001101101111010101001000101011010111000001100001110010111000110010000100011011101011000000000001000010001001001011001111111001110111111101000100001110111110110011111011100000000000001001110010011010001111101001101101000110100010110100110101010100111100111101000000101000000111010011000000110100101100110110100000001010010010011010000001100001101101100011110000010110101011000111011100111001111011010010000101110011001100000000000101001111100100110100100001100000111111000001111011101011010101101011111000010001011100111010011001000111111001101110011101110111010110000110111000100000011101100011010101000110011101101000011010110001010101111110011000101010110101010001100001011100101011100100010110011011100001010011101110001110110111001111001000111011000110000010010010101101000100010100011100111101110001001001101011010000111001101110001001110010101100100011010001111010110110000010010010010101011110000011001001110110011100000010101101011100011010100000011010110100101010110010000111011110110000011000000100111101111111010010101101001100001111010110100101100111110000101111110111111000111110111010110110001101010110111101101000001010101111010000011001101111011110000101111011000101001010101011010100000110111011000101011110001110001101000011111100101011001010110000101111100101110110101011110001111110111101100011110100010100111111011101111000101001010101110011000100111011001110001110101110011100101011101101011101101000011000100001111011100010100101010110000101100000101000000111110000011101010100001010010001111101010000110001010111100100110011100010110010011111001100011111101010000010010100001000100101010101100101100001010010101010010100110100100010111011101100011111101101101110011101010010000111101110101111110100000101010000111101110100010100010011101011010101110100110010011000110110100010101100010000010101010011101110100110011101101111000100000100001100111111001011011000001010110010111001001100100010010011100010101111011100101000111111101001011100111101111100001001001001111110110010101010111101110011000101100001111101000100101000001100111001001001110000001110111000001110110100001110111001000100001000100000001101100101001011110000111011000101110000101010101111100110011100111111010110010110011011100011111001011010111101011101001110101000110001010000010010000100001100001000010101110100111001011000110010000001010010111010011111010110000000001111110011000110000001011011111110101110101100001110100110001001011010000100100011000101011100011100010101100000101000000011011000001111010011110010001111000100100101101100010011010010000000011100111010110100000010000001000111011011101101111111011010101101010000000011001011110100101111111000111100001011010010101111001000110001111001110001001000100010001001001010111001001111111110100000111100101011011000010010001110010110111000001111011010011101111011001100111111100111000010001010101010110011011001011011010010100001110100011011100001110110101000110101011000000100101000011010011110100100101101111100000001011001111010001011110100011010011101001111100011001100001010010100001001101010001101110101011111010000011001000100110011100100011011110000111001111111101101101101111101110111110100111101110011110110101110110100010100011111011000011000100101000101100011111111010110000010100010010001010000110101011010101111010010101110010011010110000001001010000110111001111001000001110000100110001011100001011010100011101011101000001101100100010110110110011011001100011001101101110110000101001111011000111110011001111111010001000101101110111000111111001010101000011110011111001010101011100000101111101100111011001110100110111100101100101110111010010010110001101011110000111001011001100011101011011101101110000001010010001101110010000011010011100101010100100000001000110011111001101010110000011110001001010111011111110101111001101111000110111010000010001101111001000110101000111010011100000010011101010001010000010000111110011100110001101110000011111010110101101111110111001110100111000111001001010100011000001100011110001010000010010001100100001100001100101010111101101110100110110011000101110110101000000001110110011010110001110100011101101011111001101000001101111100001011110011101010000000101011101001001100001010011000101101110101010010001111110010011011011110100101111101101001000010101010100010101100010110010100001100110000011100011011111001101110110110011011000101110101010000011010000011010011000111100110001001111011001010110101100000111111111011101001111110101001011010000101011111001001001011111000001000001001110101100110011000000000010100100011000110011101110001100101010011110100110000010001100100011001001110000011100000011001111000110110100101010001001111001011001101010001100001101010100010001110110000011011001101110011101000001100001000011101111000010110111111001100010001111000011111100100010010111010000001011100111011010011110110110000110011101010001010100010110011010111000111010010100111110000110111000110000100100110001110000111110011010001010001111001100110111001011101001110101001001001011100010101001110101100000000110100110011111111110000001110101101010011001101001110100100100000000111011000110011010100010101000111000110101101011100010111011000011101010010000110011100011001011111110100000001101110100010101010101011110110001011010011001100111100110110110010100000001110110011011101100110100010000111010111011100001001001010001011000010011100011001010111101110000110001100101010111000001100010000011100100010001000111000010100110010001110110011000100110101011111011011101110001110100010101111110000100111110011110011000100001110001100110100100011011100010000000100110001000101111101010000111001001100011101110001011110010000100101101101100100001100101111001100001111010000010011010000111100001101100011000101000011100011101001101101111111001110001100011110111110100101001101101111010110101001111011111001111111101111101010101111010110111001000011000000001101111111111111101100111101010111101001000010101011010010001100010101111011111010011011110011111100101010010111110000110001010100111000101101101001110000010000001010011001011011101000111100111101100101010110001100010101101011100110000011110111111000110010011111001011111100111001011110010011010001100111111001000110110011010111010111001010000110101100101000101101110010111001110110010010011011101100010100000000001011111000001000000010100111000110101110011011100010001110101001111111010000110010101010101000010011101110101111100001000010111; 
		letterEncoding[ 5] <=10000'b1100101100111000010111110110111010011110110001110110101101001111110011101011001001111100001000011010001101011001001111101110100110001111101010110010010000110000111111111011111001011111000011101011000010011000001100000011000010101011100101110011001001000111011101000000100100111110001010101000101110100100100101000011011010000100101000111110000110100010011000011110010001001101100001111010101111111011100110001000011011110100000001100111010001111011100101101100010000111011100001111100001100011101100011010011000100000100111110111001000100011100101101011100100110111011111110110101010100111001111001000011101100110001100011000101101100011011010000101000010001101011111100100010111011011000101001111100111010000110110000001000011010101100011001111001110110011111011000011000111010101011011101000100101000110010111011010000101001000100111101111011001000100000100111100011101001011110110100000100101010011100100001101110101010011010000101101000011001100010110110000000010110100101110110000101111111100101001010111100011011011100010000011111100110110110010110101110000110011100011011011100001011101100110011011101010110000010110001011111110111110110110011101101010101111100000111100111011101011011110000010100010100101100110011000111001100111100010111000111001110111011110110101010000111111110001010000100011000101111001011011101011111010011111101110101111101110101010011101011111101010111100101010001101111000101110010011011000110100111000011111011110011100111011010110100000111111111010110110111111011001100000010100000111000011101011100000101000001110011011100100011111110010010000101101111101010101110000000100001011111100111000101100101010001110011111010110110000000101100000100001011100010101001110000111010111000110100111111011010111001101001011101110111001110001001100100000010101001101110010011000000101010010100111101111110110010110101000101101000010110000000111100010001101110110001011101100101000011100011011110001010101101100111001111101011001011011001111100100111010010001011000111011110000110000011000010010010101101110000011100110111110000100000011000101111111000001001101000001000111000000111110110011101110100011001001011000111101101111011110010110010000010010110000101111101000001000011111001010101001111111001101011110100001110011011010001010010101101100000000100100110100000011011110001101001111001000001011101010000000101011011000111100111001010011010100101100100010000010010111101100000001011111001001111111001111001001011101000001101011100000111101010001101111111010110100011000101111011100101111001001001011001110100110001011011101011111010110100001011101010100011100111100110100110100001100111001000011011000101010111110111011011001010111011101010110000100110001111110100110001001010001100010001011011110000001111110001011001011101011111100110111110111111110001110100110010011101010110100100011000100011001000101110110001010001010000011011000101101010000010111100100001010011010001111111000010011101000101101110010011010110101111101010100101100000000100100101011110001001001100101011000101010111010010010111101001010010000110010100100001110000010101110001010011010000000110001100010101100011001110111001100101011011011101001000101000010101101111101111000101001100111000000111100011010011011000000110000000000110010111001111111011000100001101010110101111000000101011000000111101100100011101101000100000010010111010010010110110000110101001001100100100111111010101101101010110000000101100001000100101101010010101011111010100001100010100001110011100010011000111000100000101111100111010011011111001011000100011100010101001010101000010111101011000000101011110010011010100011011011010000000100001000100010001101101111010101001010101011010111000001100001110010111000110010000100011001001011000000000011000010001001001011001111111101110111111101000100001110111110110011111011100000000000001001110110011010001111101011101101000110100010110100110101010100111100111101000000101000100111010001000000110100101100110110100000001010010010011010010001100001101101100011110000010110101011000111011100111001111011010010000101110011001100000100001101001111100100110100100001100000111111000001111011101011010101101011111000010001011100111110010101000111110001100110011101110111010110000111111000100000011001100011010101000110011101101000011010110001010101111110011000101010110101010001110001011100101010100100010110011011100001010011101110001110110111001111001000111011000110000110010010101101000100010100011100111111010001001001101011010000011011101110001001110010101100100011010001111110110110001010010010010101011110000011001001110110011100000010101101011100011010100000011010110100100010110010000111010010110000011001000100111101101101010010001101001101001111010110100101100111110000101111110110011000110110111010110110001101010100111101101000001010101111010000011001101111011110000101111011000101001010101011010100000110111011000100011110001010001101001011111101101011001010110000101111100101110110001011110001111110111101100011110100010100111111011101111000101001000101110011000100111011001110001111101110011110101011101101011101101100011000100001111011100110100101010110000101100000101000000111110000011101010100000010010001111101010100110001010111100100110010000010010110001111001100011111101110010010010101001000000101010101101101100001010010101010011100110100100010011011101110011111101001101110011101010010000111101110101111110100000101010000111101110100010101010011101001010101110100010010011000110110101010101000010000010001010011101110100100011101101111000100010100001100111111001011001000001010110000111001001100100010010011100010101111011100101000111111101001011100111101111100001001001001111110110010101010101101110011000101100001111101000000101000101100111001001001110000001110111000001110110100001110111001000100001000100000001101110101011011010000011011000101110000100010101111100110011100111111010110010111011011100011111001011010111001011101001110101010111001010100010000000100001100001000010101110100111001011000100000000001010110111010011111010110010010001111110011001110000001011011111010101110101100001110100110001001011110000100100011000101011100011100110101100000101000000011011000001111010001110000011111000100100101000100010011010010000000011100011010010100000010000001000101001010101101111111011110100101011000000011001001110100101111111000111100001011010010100111001000110001111001110001001000100010001001001011011001001011011110110000111110101011011000000010001110010110111000001111001010011101111011001100111111100111000010001110101010110010010001011011010010100001110100011011100001110110101000110101011000000100100000011010011010100110101101111100000001011001111010001011110101011010011101001111100010001100001010010000011001101010011101110101011111000000011001000000110011100100011011100000111001111111101101001101111101110111110100111101100011110110011110100100000100011011011000011000100001000101100011111111010110000110100001010001010000110111111010000111010010101110010011011110000001001010000110111001111011000001110000100100101011100001011010100011101011101000001101100100011110110110011011001100011001101101110110100101001111011000111110010001111111010001000101101110111000100111001010101000010110011111001010101001100000101111101100111010001110100110111100101100101110111010010010110001101011110000111001011001100011101011011101100110000101010000001101110011000011110011100101010100110000101010110011111001101010100000011110001000110111011111110101111001101111000110111010000010001101111001000110101000101000011100000010011101010001010000010110011100011100110001101111000011110010110101101011100111001110100011000011001001010100011000001100010110001010000001010001100100001000001100101010111101101110100110110011000101110110101000000001110110011111110001110000011101111011011001001000001101111100001011110011101010000000101011101000001100001010011001110101110101010010001111110010010011011110100101011101101001010010111000100010101100010110010100001000110000011100111011111001101110110110010011000101110101010000011010000011010011000111100110001001110011001010110101100000111111111011001001011100101001011010000101011111001001001011011000001000001001110101100110011000000010010100101011000110001101110001000101010011110100110001010001100100011000001110000011100000011001111000110010100001000001001111001011001101010011100001101010100010001110110000011011001001110011101000001100001000001101111000010110111111001100010001111000011111100100010010111010000001011100111011000001110010110000100111101010001010110010100011010011001111010010100111110000110111000110000000100110001110100110110011010001010001111001100110111001011101001110101001011001011100010101001110101100000000110100110101111111110000001110100101010011011101001110100100100000000111011000110011010100010101000111101110101101011100010111111000111101010010010110011010011000011011110100000011101010100010101010111011111110001011010111001100111000100110110010100000001110110011011101100110100011001111010111011101001101001010001011000010011100010001010111101010000110001110100010111000011101010000111100100010001010111000010100110010001110110011000100010101011111011011101110001110100010001111110100100111110011110011000100001110001100110100100011011100010000000101110001000101111101110000011001000100011101110001011110010000100101101101100100001100101111110100001111110000010011010000110100001101100011000101000011100001101001101101111111001110001100011110011111100101001101101101010010001001111011111001111111101111101010101111010110111001000011000000001101111110111111101100111101010111101001000010101011010000001100010001111011111010111011110011111100111010010111110000110001010100111000100101101011110000010000001010101001011011101000110100111101100001010100101100000101111011100110000001100111111000110010011111000011111100111001011110010001010001100111111001000110110011010111010111001010000110101100101000101101110010011001110110010010011011101100010100000000001011110000001000000010000111000110101110011011100010011110101001111111010000110010100010101000010011101110100111100001100010111; 
		letterEncoding[ 6] <=10000'b1100101100111000010111110110101010011110110101110110101101001111110011101011001001111100001010011010001101001001001111101110100100001111101000101010010000110000111111111011111001011111000011100011000010011000001100000011000010101011100101110011001001000101011101001000100100111110001010101001101110100100000101000011011010000000100000111111010110100010011000011110010001101100100001111010101111111011100110001000011011110100000011100111010001111011100101111100010000111011100001111101001100011101100011000111000100000100111110111001000100011100101001001100101110111011100110110101010100111001111001000111101110110001100011001100101100011011010001101100010001101011111100100010111011011000101101011100111010000110010100001001011010101100011001111001110110011101011000010001111010101011010101000100101000010010111010010000101001000100111101011011001000100000110111110011101001011110110100000100101010111101101001001111101010011010000101101000011001100011110110000000000110100101110110100101111111100111001010111100011011011100010000010111100110110110011110101110000110011100011011011100001111101101110011011101010110000110110000111111110111110110110010001101000101111100011111100111011001011011110000010100010101101110110011000111001100111100010111000111001110110011110110101011000110111110001010000000011000101101001011011101001110010011011101111100110101110101010001101011111101010111100101000001101111000101010110001011000110100111000011111011010011100111011010110100000111111110010110010101111011001100000010100000101000011101011100000101001101110011011100100011111110010010000101101111001010101110000000100001001111100111000101100100010001110111111011100110000000100100000100001011100010101001110000111010101000010100111111010010111001101001011101110111001110001001100100000010101011100111010011000000101000000000111101011110110010110101000101111000010110000000111100010001101110010001011101100101000011100011011010001010100101100101001011101011001001011011111100100110010010001011000111011110000110000011000010010011101101010000011100110111110000100010011000101111111100001001101010011000111000001111110110011101110100011001001011000111101101111011110110110010000010010111000101111101000001000011111001010001001111111001111011110100001110010011010001010010101101100000000100101110100000011011100001101000111001010000011101010000000101011011000111100110001010011010100101100100010000010010011101100000001011111001001110111001011001001011101000001101011100000111101010001101111111010110100011000101111011100101111001001001011001110100110001011011101011111010110100001011001010100011100111101110100110100001100111001000011011000111010110110111011011001110111010101010110000100110001111110101110001001010001101010011011011110000001101010001001001011100001110100100111110111111110001110100010010011100010110100100011000100011011000101111110001010001010000011011000101101010000010101100100101010011010001111111000010011101000101111110010011011110101001101010100101100000000100100101011110001001001100101011000101010111000010010111101001010010101110010000100001110100011100010001010001010000000110001101010101100011001110111001100101011011011101001000001000010101101111101111000101001110111000000110100011010011010000000110001000000110010111001111111011001100001101011010101111000100101011000000111101101100011101101000100000010010110010010010100110000110101001001100100100110111010101101101010110000001101000001000100100101011010101111111010100001100010100001110011100010011000111000100000101111100111010011011111001011000100010100000101001010101010000111101011000000101011110010011010100010010011100000000100001000100010001101101111010101001010101011010111000001100001110010111000110010000110011001001010000000010011100010001001001011001111111101110101111101000100001111111110110011111011100000000000001001110110011010001011101011101101000110100010110100110101010100111100111101000000101000100111010001000000110100101100100110100000001010010010001010010001100001001101100011110000010110101011000111001100111001101011011010010101110011001100000100001101001111100100100100100001100000111111000001111011101010010101101001101000010001011100110110010101000111110001100110001101111111010110000111011000100000011001100001010001000110010101001000011010110001010101111110010000101010110101010001100001011100101010100100010110011011100011010011101110001110110111001011001000111011000110100110010010101100000100010100011000111111010001001001101111010000011011101010001001110010101100100011010001011110110110001010010010010101011110000011001101110110110100000010101101011100011010100000011010110100100010101010000111000000110000010001000100111101100101110010001101001101001111010110100101100111110000101111110110011000110100111010110110001101000100110111101000001010001111010000111001101111010100000101111011000101001010101011100100000110111011000101101010001010001101001010111101101011001110110000101111100101110110101011110001011111111101100011110101010100110110011101111000101001010101110011000100111011001110001111101110011110101010101101011101101100011000100001111011100110100111010110000101100000101000000111110000011101010100000010010001111101010100110001010111100100110010000010010110001111001100011101101110010010010101001000000101011101101100100001010010100010110100110100100010011011101110011111011001101110011101010011010111101110101111010100000111010000111101110000010101010011101001010101110100010010011000110110101010101000010000010001010011101110100100001101111111000100010100001100111111101011001000001110110000111101001100100010010011100010101111010100101000111111101001011000111101111101001001001001111110110010101010100101110011000101100001101101000000101110101101111000001001110000001110111000001110110100001110111001000101101000100010001101110101011011010001011011000101110000101010101111100110011000111111010110010111000011100011111001111010111001011101001110101010111001010100010000000100001100001000010101110100011001011000100000000001010110111010011111010110010010001111110011001110000001011011111010101110100100001100100110001001011111000000100011011101011100011110110101100000101000000011011100001111011001110000011111000100100101000100010011010010000000011100011010010110000010010001000101001010101101111111011110100101011000000011001001110100101111101000111100001011010010100111101000110001111001110011001000100010101001001011011001001011011110110000111110101011011000000110001110010110111000001110001010011101111011001100111110110111000010001110101110100010010001011011010010100001110100001111100001110110101000110001111000000100100000010010011010100110101101101100000001011001111010001011110101011010011101001111100010001100001010010000011001101011011101110101011111000000011001000001110011100000011011100000111001110111101101001101101001110110110100111101100011110110011110100100000101011011011000011100100001000101100011111111010110000110101001010001010100110111111010000101010010101110010011011110000001001000000110111001111111000111110000100100101111100001011010100011101011101000001101100100011110010110011011011100011001101101110110100101001111011000111110010001011110010001000000101100111000100111001010101000010110011011001011101101100001101111111100111010001110100110111000101100101110111010010010110001101010110010111001011001100011101001011101100110000101010000001101110011000011110011100101010100110000101010100011111001101010100000011110011000100111011111110101111001100111000110111010000010001101111001000110111010100000011100000010011101010001010000000110011100011110110001101111000111110010110101101011100111001110100011000011001001010101001000001100010110001010000001010001101100001000001100100010111101101110100100110011000101110100101000000001110100011111111001010000011101111001001001001000001101111101001011110011101010000000101111101000001000001010011001110111110101010010001011110010010011011110100101011101101001010010111000100010101100000110010101001000110010011100111011111001101110110110010011000100110101000000011010000011010011000111100110000001110011001010110101100000111111111011001011011100101011011010100101011111001011001011011000101000001001110101110110010000000010010100101001000110001101110001000101010011110100110001110001100100011000001110000111100000011001111000100010000001110001001111001011001101000011100001101010100010001110110000011011001001110011101000101100001000001101111000010110111111001100010001111000011111100100010010111010000001011100111001000001110010110000100111101010001010110010100010010011001111010010100111010000010111000010000000100110001110100110110011010001010001110101110111111001011101111110101001011001011100010101011110101100000000110100110101111111110000001111100001010011011101101110000101100000001111011000110011011100010101000111101111101101011100010111111010111111010010110110011010011000011011110100000011100010100010101010111111111110001011010111001110111000100110110010100000101110110011011101100110100011001111010111011100001101001010001011000010011100010001010111101010000110001110100010111010000101010000111100100010001000011001010100110010000110010011000100010101010111011011101110010110100010000111110101100111110010110011000100001110001100110100100011011101010000000101110001000101111101110001011001000100011101110001011110010000100101101101100100001100101111110100001111110000010011010000110100011101100011000101000111000001101001101001111111001111001100011110011111100100000101101101010010000000111011111001111011101111101010101111010110101101000011000000001101111110111110101100111101010111101001011010100011010000001100010001111011111010011011110011111101011010010101110000110001010100111000100101100001110000010001011010101001011011100000110100111101100001010100101000000101111011100110000001110110111000110010010111000011111100111001011110010001010001100111111001000110110011010111010111001010000100101100101000101101110010010000110110010010011011101100010100000000001011010000101000000010000111000110101110011011100010011110101001111111010000110010100010101000010011101110100111100001100010110; 
		letterEncoding[ 7] <=10000'b1100001100111000010111110110101010011010110101110110111101001111100011101011101001111100001010011010001101001001001111101110100100001111101001000010010000110000111111111011110001011110000010100011000010011000001100000001000010001001100101110011001001000101111101001000000100011111001000100001101110100100000101000010011010001000100000111111010110110010011000011110010001101100100001111010101111011010100110001000011011110100000011110111010001111011100101111100010000111011100011111101001100011101100011000111000100000100101110111001000100011100101001001100111110111011100110110101010100111001110001000111101110110001100011001100111100111011010011100100010001101011011100100011111011011000101100001100111010000110010100001001011010101000011001111001110111001101011001010001101010001011010101000100101000010010111010010001101001000000111101011011001000100000010111110011101001001010100101000100101010111101111001001111101010011010000101101011011001100011110110000001000110100101110110000101111111100111001010111100011011011100010000010111100110110010011110101110000110011100011011011100001111101101010011010101010110100110110000111110110111110110110010001101000101111100011110100011011001011111110000010100011101101110110011000111001100111100010111000111001110110001110110111011000110111111001010000000011000100101001011011101001111010011011101111100110101110101010001101011111101011111100101000001111111000101110110001011000110100011010011111011010001100111011010110100000111111110010110010101111011001100000010100001001000010101011100100101001101010011011100100011111110110010000101101101000011100100000000100001001110100111001101100100010001111111111011000010000010100100000100011011100010101001010000101010101000000100111111011000101011101001011000010111001110001001100100000010101011101111010011000000100000001010111101011110110000110001000101111000010110000000111100010001001110010001011101100101000011100011111010001010100001100101001011101011001101001011110100100110010010001011000111001110000110000011000010010011100101010000011000110111110000100110011000101111111100001001101010001100111000101111110100011101110100011001001011000111101101111011000110110010000010010111000101111101000001000011111001110000101111111001111011111100001110010011010001110010101101100010000101100110100000011011100001111000111001010000011101010000000101010011000111100110001010011010100101100111010000010010011100100000001011111001001110111001011001011011101000001101011100000111101010001101111111010111100011000100111111100101111001001001010001110100110001011011101011101010010100001011001010100011110111101110100110100001100111001001011011001111010110110111011010001110111011101010110000100110001111110101110001101010001101010011011001110000001101010001011000010100001110100100111110111111110001110110010011011100010111100100011000100011011000100111110001010001010000011011000101101010000010101100101101010011010001110111000000011101000101111100010111011110101000101010100101110000100000100101011110101001001100111011000101110111001010010101101001010010101111010000100001110100011100010001011001010000010110001110010101100011001110111001100101011001011101001000001000010001101111101111000111001110111001000110100011110011010001000110001000000110010111001111111111001100101001011010101111000100101011000000111101101100011101101000100000010001110010000010100110010110101001001100100100110111010101101101010100000001101000001000110110101011010101111111010100001100010100001100011110010011010011000100000101111000111010011010111001011000100010100000101001010101010000111101011010001101011110010011010100010010011100000000100001000101110001111101111110101001010101011000111000001100001110010111000110010000110011001001010000000110011100010001001001010101111111101110101001001000100001011111110110011111011100000000000001001110110011011001011101011101101000110100010110101110101010100111100111101000000100000000111010001000000110100101100100010100010001010010010001011010001101001001101100011100000001110101010000111101100111001111011011011010101110011001100000100101101001111100100110100100001101000111111000101110011101010010101101001101000010001011100110010010101100111110001100110001101111111010110000111011000100000011001100001010001000111001101101000011010110001110111111110010000101010110101010001100001011100101010100100010110011011100111010011001110001110110111001011001000111011000110100110010010100101000101011100011000111111010001001001101011000000011011101110001001110010001100100011010001010110110110001010000010010111011110000011001101110110110100000010101101011100011000100000111011110100100011101010000111000001110000010001000100111101100001100010001101001101001111010111100101101111110000101111111110011000110100111010110110001001000100111111101000001010001111010110111001101111010100100111111011000101001010101011100100000110111011000101001110001010001101000010111101101011001110110000101111100101110110101011110001011111111101100011010101010100110110011101111010101011010101110011000100111011001110001111101110011110101000101101011101101100011000100001111011110110000110010110000000000000101000000111010000011101010100000010010001111101010100110001011111100000110010000010010100001110001100011101101110010010010101101000001101011101101100100000111010100110110100110100101010011011101110011111011001111110011101010011000111101110101111110100001111010001111101110000010101010011101001110101111100110011011000111110111010101000110000010001010111100111100100001101111111000100010100001101111111100011001000001110110010111101001100100010010011100010101111010100101000111111101001001000111101111101001001101001111110100010101010100100110011000101100001001001000100101110101101111000001001110000001110111000001110110100001110111000000101101000100010001101110101011011010001111011000101010000101011101111100100011100111110010110010111000011100011110001111010111001011101001110101010110001010100010000100100001000001000010101111100011001011000100001000001010110011010011111011110000010001111110011001110000001011011111010101110100101001100100110001001011111000000100011011101011100011110110101100000101000100011011100001111111001010000011101000100100101000100000011011010000000011100011010000111000010000001000101001010101101111111011110000101011000000011001001110100100111101000111100001011010010100101001000110001111001110001001000100010101001001011011001001011011110110000101110101011011000000110001110011110111000001110001010011101111011001100111101110111000010001110101010100010010101011011010010100101110100001101100001110110101000111001111000000100100000010010011010100110101101101100000000011001101010001011110101011110011101001111100110001100001010010000010001101011011101110101011111100000011001000001111011100000011011000000111001010111101101001001101001110110110100111101100011110110011110100100000101011011011000011100100001000101100011111111010110000110101001010001010100110111111110000101011010101110010011011110000001001010000110111001111111000101110000100100101111100001011010100011101011101000001101100100011110010110011011011100011001101101110110101101001111001000111110010001011110010001000000111100011000100010101010101000010110011011001011101100100001101111111100111010001111100110111000101100101110111010010010110001111011110010101001011001100011101001011101100110000001011001001100110011000011110011100101010100110100101010100011110001101010100000011110011000100111011111110101111001100101000110111010000010001101110001000110101010100000011100000010011101110001010001000110011100011110110001101111001111100010110101101011100111001110100011000011001001010101001000001100010110001010000101010001101100001000001100100010101101101010100100110011000101110110101000000001110100011111111001010000011101111001001001001000001001111101000011110011101010000010101111101000001000001010011001110111110101010010001011110010010011011110100101011101101001010010111001100010101110000110010101001001110010011110111001111001101110110110010011000100110101000000011010010011010011000111100110000001110011001010110111100000111111111011001011011100101011010010100101011111011011001011011010101000001001110101110110010000000010010100111001000110001101110000000101010011100101110001110011100100011000001110010111100000011001111000100010010001100001001111001011001101000011100000101010000010001110110000011011001001110011101000101100101000101101111000010110111111001100010000111000011111100100010010111010000101011100111001000001110010110000100111101010001010111010100010010011001111010010000111000000010111000010000000000110001110100110110011010001010001110101110111111001011101110110101000011001011100010111011110101100000000100100110101111111110000001111100001110011011101101110000101100000001110011000110011011100010101000111101101101101011100000011111010111111010010110110011010011000011011110100000011100010100010101010111110111110001011010111001110111000100110110010100000100010110011011101100110100011001111010111011100001101010010101011001010011100010001000111101010000110001010100010111010000100000000111100100010001100010001010100110010000110010011000100010101010111011011101110010110100010000111110101100111110010110011000100001110001100110100001011011101010000000101110101000111111101110001011001000100011101110000011110010110100101001101100100001100101111110100001111110000010011010000010100011101100001000101000111100001101001001001111101001111001100011110011111100100000101101001010010000000111011111001111011101111101010101110111110101101001011100000001101111110111110101100111101010111111001011010100011010001001100010000111011111110011011110011111111011010010101110000010001010100111000100101100001110000010001010010101001011011101000110100111101000011010000101000000101111011100110000001110110111000110010011111000011111100111001011110010001010001100111111001000110110011010111010111001010000100101100101001101101110010010000111110010110011001101100010100000000001011010000101000000011000111001110101110111011100010011110101000111110010000010010100010101001010011101110100111100001100010110; 
		letterEncoding[ 8] <=10000'b1100001100111000010111110101101010011010110101110110111101001101100001101011101001111100001010011010001101001001000110101110100100001111101001000000010000110000111101111011110001010110000010100011000010011000001110000001000010001100100101110011001001000101111111001000000110011111001000100001101110000100000101001010011010001000100000111111000110110010011001011110010001101100100001111010101111011010100110001000011011110100000011110111010001111011000101111100010100111011100011111101001100011101100101000111000101000100101110111001000101011100101001001110111110111011100110110101010100101101110001000111101110110001101011001100111101111001000011100100010001101011111000100011011011011100101100001100111010000110010100001001011011101100011001111001111111000001011001010001101010001011011101000100101000010010111010010001101101010000111101011011001000100000010111110011101001001010100101000100101010111101111001001111101010011110010101101011011001100011110110000001000110100101110110000100111101100111001010111111011011011100010000010111100110110010011110101110000110011100011011011100001111111101010111010101010100100110110010011110110110110110110010001101000101111000001110100111001001011111110000010100011101101110110001000111001100111100010111000111001110110001110100111011000100101111001010000100011000100101001011011101001111010011011001111100110101110111010001101111111101011111100100010001111011000101100110001010100110100011010011111011011001100111011000110110000111111110010110011101111010001100000010100001001000010101011100100001001101010011011100100011101111110010000101101100000001100000001000100001000100100111001101100100010000111111111011000010000010100100000100011011100010101001010000111010111001000000111111011000101011101001011000010111001110001001100100000010101011101111010011000000111000001010111101011110110000110001000101111000010110000010111100011001001110010001011101100101000011110011111001001001100001100101001011001011001101001011110100100100010010001011001111001110000110000001000010000011100111010000011000110111110000100110011100101111111100001001101010000100111000101111110100011101110100011011001011000111101100111011000100110010000011010111000101111101000000000011111001110000101111111001111011111100011110010011110001110010101001100010000101100110100000011011100001111000111001010000011101010000000101010011000111001110001010011010100101100111010100010010011100100000001011111001001110111001011000011011101000001100111110000111101010001101111111010111100011001100111111100001011001001001010001110100110001011011101011101010010100001011001010100011110111101010100010100001101111001001011011001111010110110111011010001110111011101010110000100110001111110101110000001010001101010011011001110000001101010011011000110100001110100100101110111101110011110110010011011100010111100100011000100011011000100111110001010001010000011001000101101010000010101100101101010011010101110111000000011101000101111100010111011110101000101010000101110001100000100101011110101001001110111011000101110111001110010101101001010010001111000000100001110100011100010001011001010000010111001100010101101011001110111000100111011001011101001000001000010001101011101111000111001110111001000110100011100011010001000010001000010110010111000111111111001100101011011010101101000101101011001000010101101100001101101000100000010011110010000010100110010110101001001100100100110110010101101101010100000101101000001001110110101011010101111111010110011100000100001101011110010001000011000100000101111000111010011010111001011000100000100000101001000101010000111100011010001111011110110010010100010010011100000000100001000101110001111001111110111001000101011000111000001100001100010111000100011000110011001001000000000110011100010001001001010101111111111110001001001000100001011111110010011111011100000000000001001110110011011001010101011101001000110100010111101110101010100111100111101000001110000000111010001000000100100101101100010100110001010010010001011010001001001001101100010100000001110101010000111101100111001111011011011110101110011001100000100101101001111110101110100101001101000111111000101110011101010010101101001101000010001011100110010010101100111110001100110001101111111010110000111011000100000011001100001010001010111001101101000011010110001110111111110110000101010110101010101100001111110001011110100010110011011100111010011001110001110110111001011101000111011000110100110001010100101000101011100011000111111010001000000101011000001011011101110001001010010001100100011110001010110110110011010000010010111011110000011011101110110111100000010101101011100011000100000111011110100100011101010000011000001110000010001000100111101100001100010001001001101001011010111100101101111111000100111111110010000110100110010110110000001000100111111101000001010001111010100111001101111010100100111111001000100001010101011100100001110011011000101001110001010001101000010111101101011001110110000101111100101010110101011110001011110111101101001010101000100110110011101111010101011010101110011000000111011001110011111100110111110101000101101011101101100011000100001111011010110000110010111000000000000101000100111010000011101010100000110010001111101010100010001011111101000100010000010010100001110001100011101101110010010010101101100001101011101111101100000111010100110011000110110001010011001101110011101011001111110011101010011000101101110101100110100001111010001111101110000010101010011101001111101111100110011011000111110111010001000010000010001010111100111100110001101111111000100010100001101011111100011001000001110110010111101001101100010010011100010101111010101101000111111101001000001111111111101101101101000111110100010001010100100110011000111100001000101000100101110001101111000001001110010001110111000001110110100001110110000000101101000100010001101100101011011010001111011000101010000101011101101100100011000111110010110010111000011100011110001110010111001011101000110111010110001010100010000100110001101101000010101111100011001011000100001000001010100111110011101011110000010001111110111001110000001011010110010101110100101001100100110001001011111000000100011011101011100011110110101100000101000000011011100001101111001000000011101000100100100000100000011011010000000010100011010000111001010000001010101001010101101111111111110000101011000000011001001010100100100101000111100001011010010100101001000110001111001110001001000110010101001010011011100001011011110110000101110101011011000000110001110011110111010001110001110111101111001001110111100110111000000001100101010100010011101011011010010100101110100001101010001110110101000111001111000000100100000010010011010100110101101101100000000011001100010001011110101011110011101011111000110001110001010011000010001101011011101110101111111100000011001000001111011100001011011000000111000010111101101001101101011110110110100111101100011110110011110110100000100011011011000011100100001000101100011111111010111000110101001010001010110110111111110000101011010101110010111011110000001001010000110101001111111000101010000100100101111100001010110000011101001101000101101100100011110010110011010011000011001101101110110101101001111001000111110011101011110010001000000111100011000100010101010101000010110011011101011101100100101101111111100111010001111100110111000101100101110111010010010110001111011111010101001011001100001101001011101100110000001011001001100100011000011110010100101010101110100111010100011110001101010100000011110001010100111001111110101111001100101000110110010000010000100110001010110101010100000011100001010011101110001010001000110001100011110110001101101001111100010110101101011000110001110000011000011011001010101001000001100010110001010000011000001101100001000001100100011100101101010100100110011001101110110101000000001110100011111111001010000011101111001101001001000000001101101000011110011101010000010101111000000001000001010011001110111110101010010001011110010010011010110100101011101101001010010111001100010101110010100010101001001110010011100111101111001101110110110000011000000110101000000111000010011010011100111100110000001110011001110010111100000111011111011001011011100101011010010000101011111011011001011011010101000001001110101110110000010000010010100111101000110001101110000000101010001100101110001110011100100011000001110010111000001011001111000100010010001100001001011000010001100000011100000101010000000001110110000011011001001110011101000101100101100101101110000010110111011001100010001101000011111100100010010111010000101111100111001000101110010110010100111101010001010111010100010000011001111010010000111000000010111000010001000000110001110100110110011010001010001110101111111111100011101110110101001110001011100010101011110101100000110100110110101111111110000001111100001110011011011101100000101100000001110011000110001011100010001000111101100101101011100000011111010111111010000110110011010011000011011110100000011100010100010101010111110110110001011010101001110111000100010110010100000100000010011011101100110100011001111010111011100001101011010101010001010001100010001000111101010000110001010100010111010000100000000111000100010001100010001010100110010000110010011000100010110010111011011101110010110100010000111110101100011110011111011000100001110001100110100001111011101010000000101110101001111011101110011011001000100011101110000001110010110100101001111100100001100101111100100001111110000010011010000110100011101100001000101000110101001101001001001111001001110001100011110011111100100101101101000010010000000101011111001111011101111101010101110011100101101001011100010011101111110111011101100111101001111111001010010100011010101001100010000111111110110011011110011111011011010010101110000010001010101111000100101100001110000010001010010101001011010101010110100111100000011010100101100000101111011101110100001110110111000110010011101000011111100111001011110010001010001100111111001000111110011010111011111001010000100101100101001101101110010011000111110010110011001101100010100001000001011010000101100000011010111001110101110111011100010011110101000111110010100010010100010111001010010101111100111100001100010110; 
		letterEncoding[ 9] <=10000'b0100001100111000110111110101101010011010110100110110101101101101100001101011101000111100001010011010001101000000000110101110100100001111101001100000000000110000111111111011110001010110000010100011000010011000011110000101000010001000100101110010001001000101111111101000000110001111001000100001101110000100000001001010111010001010100000110111000110110010011001011110010001101100100001111010001111011010100110001000001011100100000010110111010001111011000101111100010100111011100001011101001100011101100101000111000101000100001110111001000101011100101001001110111110111011100110110101010100101111110001001111101110110000001011001100111101111001000011100100010001101011111000100011011101111100101100001100111110000110010100001001011011101100011001111001111110000001011001010001101010001011011101000100101000010010111110010001101101010000111101011010001000100000010111100011101011001010110101000000101011111101111000001111101010011110010101101011011001100011110100000001000111100101110110000000111101100111001000010111011011011100010000010111100110110010111111101110000111011101011001010100001111111101010110010101010000100110110000011110110110110110110110001101000101111000001110100111001001011111101000010100011101101110010001000111001100110100010111000111001010110001110000111011000000101111001110000100011000100001001011011001001110010011011001111100110101110111010001100111111101011111100000010011111011000101100110011010100110100011010011111011011001100111011000110110000111111110010010101101111010101100000010100001001000010101011100110001001101010011010100100011101111110110000101101100000000100010001000100001000100100111011101100100010000111111111010000110000010100100000100011011100010101001010000101010111001000000111111011000101011101001011010010111001110001001100100000010111011101111010011000000111000000010111101011110110010110001000101111001011110000010111110011001001110110001001101100101001011010011111001001001100001100101001011001011001101001010110110100100010010001011011111001110000110000001001010000011100111010010011100110111110000100110011100101101111100011001101010000100111000101111110100011101110100011011001011000111101101111011000100110010000011010101000101111101001000000011111001110000101101111001111011111100011110010011110001110010101101100010000101100110100000010011101011111000111001010000011101010000000101010001000111001110001000011010100101100111010100011010011110110000011011111001001110111001011000011011101000001100101110000111101010001101111111010111100011001100111111100001011001001001010001110100110001111011101011100010010100001011010010100011110110101010100010100001101111001101011011001111010110000110011011001110111011101011110010100110001111110101110000001110001101011011011001110000001101010111011000110100001110100100101110111001110011110110010011011100010110100100011000100011011000100101110001011001010010011001001101101010000010101100101100010011010101110111000000001101000101111100010110011110101010100010000101110001101000100101011110101001101110111011000101110111001110010101101001110010001111000000100001110100110100000001011001000100010011001100010001111011001110101000100111011001011101001000001000010101101011101111010111001110111000000110110011100011010001000010001000010110010111000111111111001100101011011010101101100101101001001000010001101100001101101000100000010011010010000010000110010110101001001100110100110110011101101101010100000101101000001001111110101011010101111111000110011100100100001110001100010001000010000100000101111000111010001010111001011000100000100000101001000100010000111000111011101111011110110010010100010010010100000000000000010101100001111001111110111011010101111000011000001100001100010111000000011000110011001000000000000110110110010001001001010101111011111110001001001000100001111111110010011111011100000000000001001110110011011001010101011101001000110000010101101110101010100111100111101000001110000000111000001000000100110101101100010100110001010010010011011010001001001001101100110100001001111111010000111101100111001111011011011110101110011001101000100111101001111110101110100101001101000111111000101110011101011010101101001101000010001011100110010111101100111110001100110001101110101010110000111011000100000011001100001010001011111001001110000011000110001110111111110110000101011110101000101100101101100001011110100010110011011100111010011001110001110110111001011101000111010000110100110001010100101000101011100011000111111010001000000101011000001011011001110001001010010001100100011110001010110110110011010000010010111111010000011011001110110111100000010101101001100011000100000111011110100100011101010000011010001100000010001000100111101101001100010001011001101001011010111100100101111011000100111110110010000110100110010110110100001000100111110101001101010001111010100111001101111010100100111111001000100001010101011100000001110011011000100001110001010001101000010111101101111001110111000101111100101010110101011110011011110111101101001010101000100110100001101110010101011010101110011001010111011001110011111100110100110101000101101011101101100011000100000111011010110000110010111010000000000101000100111010000010101010100000111010001101001010100010001011111101000100010000010000100001110001100011101101110010010010101101100001100011101111101100000111010100110011000110010001010011001101110011101011001111110010101010011000101001110101000110100001111010001111100110000010101010011101001111001111100010011011000111010111010001010010000010011010111100111100111001101111111000100010100001111011111100011001000001110110010111110001101100010010011100010101111010101101001111111101001000001111111111101101101101000111110100010001010100100110011000111100001000101000100101110001101111000001001111010001110101000001110110100001110110000000101101000100010001101100101011011110000111011011101010000101011100001100100010000111110010110010111000011100001110001110010111001011001000110111010110000010100010000100110001101101000010101111100011001011000100001000001010110111110111101011110000010001111110111001110000001011000110010101110100101001100100110001001011111000000100011011101011100011110110101100000101000000011011100001001111101000000011101000100100000000100000011011010000010000100011010000111001010000001010111000010101101111111111010000101011000000011001001010100100100101000111101001111010010100101001000110001111001110001001000100010101001010010011100001011011110111000101110101011011000100111001110011110111010001110001110011101111011001110111100110011000000001100101010100010011101011011010011100101110100001101010001110110101000111001111000000100100010010010010010100110101101101100000000001001110010001011110001011110011101011111001111001111001010011100010001101011011101100100011111100000011001000001101011100011011011000000111000010101101101001100101011110110110100111101100011110110011110010100000100011011011000011101101001000100000011111111010111001110100001010001010110111101111110000001011010101110010111111110000000001010000110101001111111000101010000100100101111100011010110000011101001101000101101100000001100000110011010011000011001101101110110101101001111001000111110111101011110010001000000111100011000100011101010101000010110011011101011101100100101101111101100111010001111100110010010101000101110111010010010110001111011111010100001011001100001101001001101100110001001011011001100000011000011110010100101011101110110111010100011110001101010100000111110000010100111001011110101111001100101000110110010000110000100010001010110101010100000011100101010011101110001010011000110001100011110110001101101010111100010110101101010000110001110000011001001011001010101001100001101010110000010000011000001001100001000001100100111100101101010100100110011001101110111101000000001110000011111111001010001011101111001101001001000100001111101000011110111010010000110101111000000001000001010011010110111110101010010001011110010010011110111100101011101101001010011111001100110101110010100000100001001110010011100111101111001101110110110000011000000110101000000111000010011010011100111100110000001100011001110000111100000111011111011001011011100101011010010100101011111011011000110011010101000000001110111110110001010000010010100111101000110001101100000100101010001100101110001110011100100011000001110010111000001011001111010110010010001100001001011000011001100000011100000101010000000001110110000011011001001110011101000101100101100101101110000010110111011001100010001100001011111100100010010111010000101111101100011000101110010110010100111101010011010101010110010000001011111010010000111000000010111000010001000000110001110100110110011010001010001110101111111011100010101110111101001110001110100010001011110101100000110100110111101111111110000001111100001111011011011101100000101100000001110011000110001011000010001000111100000101101011101001001111010110011010010110110011010011000011011110100000011100010100010101010111110110110001011010101001010111000100010110010100100100000010011011101100100100011001111010011010100001101011010101010000110001100010001010111100010000010001010100000111010000100000000111000100010001110010000010100110010000110010011000100010110010111011011101110010110100010001111110101100011110011011011000101001110001000110110001111111101010000000101110101001111011101110011011011000100111101010001001110010110100101000111100100011100001111100110001111110000110001010000110100011101100101000100000110101001101001001001111001001110001100011110011111100100101101101000010010000000101010111001111011101111101010101110011100101101011011100010111101111110111011101100111101001111111001010010100011010101001100010000111111110110011011110011111011011010010101110001010000010101111000100101100001010000010001110011111001011010101010000100111100100011010100101100000101111011101110110001110110111000110000011100000011111100111001000110010001010111100011111001000111100011000111011111001010000100101100101001101101110010010000111110010110011001001000010100001000001011010000101100000011010111001110101110101010100010011110100000111110010100010010100010111001010010101111000111100001000110110; 
		
	end 
end


always @(posedge clk) begin
	if (rst) begin
		letterVector <= letterEncoding [inputLetter];
	end
end
 
endmodule
